* PEX produced on Sun Apr 16 07:15:33 PM CEST 2023 using /foss/tools/iic-osic/iic-pex.sh with m=1 and s=1
* NGSPICE file created from hpretl_tt03_temperature_sensor.ext - technology: sky130A

.subckt hpretl_tt03_temperature_sensor io_in[1] io_in[2] io_in[3] io_in[4] io_in[5]
+ io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6]
+ io_out[7] io_in[0] vccd1 vssd1
X0 temp1.capload\[7\].cap.Z temp1.dcdc.Z a_6736_15055# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X3 vssd1 a_1766_2223# clkbuf_1_1__f_io_in[0].A vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X7 vccd1 a_2198_1653# a_2125_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X11 a_3312_18793# a_3063_18543# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X29 vssd1 io_in[0] a_1766_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X30 a_3656_20407# temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref.TE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X32 _095_.CLK a_1674_1135# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X48 a_4130_1653# a_3971_1679# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X53 a_3404_17999# a_3155_17999# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X54 temp1.capload\[2\].cap.Z temp1.dcdc.Z a_8004_16617# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X57 a_2125_1679# a_1591_1685# a_2030_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X65 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref.Z temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[4\].pupd.A a_3312_18793# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X67 vccd1 a_1766_2223# clkbuf_1_1__f_io_in[0].A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X71 vssd1 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[4\].pupd.TE a_3331_19407# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.235625 ps=1.375 w=0.65 l=0.15
X81 a_2321_10703# _055_.A1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X92 _051_.Y _051_.B1 a_3615_21263# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X93 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref.Z temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[4\].pupd.A a_3240_17455# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X100 a_5796_16911# a_5547_16911# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X104 a_4337_1135# _061_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X107 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref.Z temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[4\].pupd.A a_3404_17999# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X111 vssd1 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref.TE a_1867_17455# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X112 vssd1 _109_.A temp1.dac.parallel_cells\[1\].vdac_batch.einvp_batch\[1\].vref.TE vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X117 _090_.A1 a_4776_14165# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10025 ps=0.985 w=0.65 l=0.15
X123 a_4535_14735# _080_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1475 ps=1.295 w=1 l=0.15
X129 vccd1 a_1674_1135# _095_.CLK vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X130 vssd1 clkbuf_1_1__f_io_in[0].A a_1674_1135# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X131 _066_.A_N _046_.A a_4413_20719# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X135 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref.Z temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref.Z a_2044_17455# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
R0 vssd1 temp1.capload\[8\].cap.TE sky130_fd_pr__res_generic_po w=0.48 l=0.045
X144 _093_.CLK a_1674_2767# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X147 vccd1 a_2956_11445# a_2890_11471# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.165 ps=1.33 w=1 l=0.15
X148 a_1840_16911# a_1591_16911# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X156 vssd1 a_1674_2767# _093_.CLK vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X158 a_4417_13353# _071_.C a_4345_13353# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.0441 ps=0.63 w=0.42 l=0.15
X160 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref.Z temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref.Z a_5796_16911# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X168 a_5072_14441# _071_.C a_4988_14441# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X170 clkbuf_1_1__f_io_in[0].A a_1766_2223# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X173 vssd1 temp1.dac.parallel_cells\[1\].vdac_batch.einvp_batch\[1\].vref.TE a_5547_16911# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
R1 vssd1 temp1.capload\[7\].cap.TE sky130_fd_pr__res_generic_po w=0.48 l=0.045
X175 a_1644_21781# _110_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X176 a_1860_16367# temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref.TE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X178 vssd1 _048_.A _112_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X182 vccd1 a_2835_25236# _114_.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X188 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref.Z temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref.Z a_1840_16911# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X200 vccd1 a_4558_1653# a_4471_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1218 pd=1.42 as=0.09135 ps=0.855 w=0.42 l=0.15
X204 vssd1 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref.TE a_1591_16911# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X210 vssd1 _080_.A2 a_2300_15095# vssd1 sky130_fd_pr__nfet_01v8 ad=0.122275 pd=1.08 as=0.05355 ps=0.675 w=0.42 l=0.15
X227 vccd1 a_1674_2767# _093_.CLK vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X243 a_2779_20175# temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref.Z temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref.Z vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.27 ps=2.54 w=1 l=0.15
X245 temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[1\].pupd.A _083_.C_N a_3345_13353# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X251 vssd1 io_in[7] a_1591_13647# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X269 io_out[6] a_2840_26677# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X272 a_3380_19319# temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[4\].pupd.TE vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.32075 ps=1.685 w=0.42 l=0.15
X276 vssd1 _090_.A2 a_4418_16367# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X277 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref.Z temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref.Z a_7656_14191# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X278 a_3421_12559# input7.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1525 pd=1.305 as=0.26 ps=2.52 w=1 l=0.15
X294 _044_.A a_2327_21807# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X298 vccd1 _085_.A1 a_4443_15529# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X302 _065_.A a_2139_10205# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X304 del1.delay_chain\[0\].inv2.A _111_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X307 vssd1 _066_.A_N a_2095_22657# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X310 a_2777_14237# _109_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.10785 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X315 vssd1 temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[3\].vref.TE a_5547_16367# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X320 a_2103_11989# _048_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.3275 ps=1.655 w=1 l=0.15
X321 a_2187_10901# _061_.B1_N vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0714 ps=0.76 w=0.42 l=0.15
X326 vssd1 a_1674_1135# _095_.CLK vssd1 sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X328 vccd1 a_1920_28853# io_out[7] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X334 _071_.C a_3512_12559# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X339 a_2927_11092# io_in[5] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X344 vssd1 _051_.B1 a_2229_9839# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X347 vccd1 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[4\].pupd.TE a_3063_18543# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X353 clkbuf_1_1__f_io_in[0].A a_1766_2223# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X364 vccd1 _051_.B1 a_5353_12265# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X367 a_3607_20175# temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref.Z temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref.Z vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.27 ps=2.54 w=1 l=0.15
X370 a_5323_17973# _092_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.1625 ps=1.325 w=1 l=0.15
X372 vccd1 del2.delay_chain\[1\].inv2.Y del2.delay_chain\[2\].inv2.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X374 clkbuf_1_1__f_io_in[0].A a_1766_2223# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X375 vssd1 _110_.A a_3065_12021# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X384 _046_.A del2.delay_chain\[3\].inv2.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.25
X389 del2.delay_chain\[0\].inv1.A a_2879_9839# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X395 vssd1 _090_.A2 a_2852_16373# vssd1 sky130_fd_pr__nfet_01v8 ad=0.122275 pd=1.08 as=0.05355 ps=0.675 w=0.42 l=0.15
X400 _093_.CLK a_1674_2767# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X403 vccd1 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[4\].pupd.TE a_3063_17455# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X407 io_out[0] a_2932_21237# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X420 del2.delay_chain\[3\].inv2.A del2.delay_chain\[2\].inv2.Y vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X421 vssd1 temp1.dac.parallel_cells\[0\].vdac_batch.einvp_batch\[0\].pupd.TE a_7931_13967# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.235625 ps=1.375 w=0.65 l=0.15
X423 a_1674_2767# clkbuf_1_1__f_io_in[0].A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X426 vccd1 _085_.A2 a_2233_15939# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.074375 ps=0.815 w=0.42 l=0.15
X431 vssd1 a_2007_11690# _063_.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X434 a_4931_1501# a_4149_1135# a_4847_1501# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X436 a_9384_16617# a_9135_16367# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X437 _076_.X a_2877_14455# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.122275 ps=1.08 w=0.65 l=0.15
R2 temp1.capload\[9\].cap.TE vssd1 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X440 a_1757_3311# a_1591_3311# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X444 a_2927_11092# io_in[5] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X463 _095_.CLK a_1674_1135# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X470 vssd1 _069_.A a_2879_9839# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X483 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref.Z temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref.Z a_9384_16617# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X489 vccd1 _051_.B1 a_2987_14735# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X491 a_8004_16617# a_7755_16367# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X494 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref.TE _090_.A1 a_4418_16367# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X495 _111_.A a_4558_1653# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.092625 ps=0.935 w=0.65 l=0.15
X496 vssd1 del2.delay_chain\[0\].inv2.A del2.delay_chain\[1\].inv1.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
R3 temp1.capload\[2\].cap.TE vssd1 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X507 vssd1 a_2835_25236# _114_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X516 a_7564_18319# temp1.capload\[9\].cap.TE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X517 vssd1 temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[3\].vref.TE a_2963_17231# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.235625 ps=1.375 w=0.65 l=0.15
X519 io_out[5] a_2104_26677# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X540 vccd1 a_1674_1135# _095_.CLK vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X544 a_3204_13879# _079_.C vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X547 _093_.CLK a_1674_2767# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X559 a_4784_17705# a_4535_17455# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X565 a_4445_11587# _071_.C a_4350_11587# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.06825 ps=0.745 w=0.42 l=0.15
X573 a_2455_1679# a_1591_1685# a_2198_1653# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X574 clkbuf_1_1__f_io_in[0].A a_1766_2223# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X575 a_2581_3311# a_1591_3311# a_2455_3677# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X589 vssd1 a_2198_1653# a_2156_2057# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X596 _048_.B a_3983_18543# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X599 a_2238_13763# _060_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X601 vccd1 _095_.CLK a_3983_1135# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X607 clkbuf_1_1__f_io_in[0].A a_1766_2223# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X611 vccd1 a_3983_18543# _048_.B vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1425 pd=1.285 as=0.135 ps=1.27 w=1 l=0.15
X612 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref.Z temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[1\].pupd.A a_4784_17705# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X616 _081_.X a_2141_14851# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.122275 ps=1.08 w=0.65 l=0.15
X618 vssd1 a_1766_2223# clkbuf_1_1__f_io_in[0].A vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X627 vssd1 _046_.B _113_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X628 a_8299_18319# temp1.dcdc.Z temp1.capload\[1\].cap.Z vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.1755 ps=1.84 w=0.65 l=0.15
X631 vssd1 a_4215_11703# _075_.A1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.17875 ps=1.85 w=0.65 l=0.15
X641 vccd1 a_1674_2767# _093_.CLK vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X651 a_2198_3423# a_2030_3677# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X654 a_2932_21237# _109_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X655 vssd1 _109_.A temp1.dac.vdac_single.einvp_batch\[0\].pupd.TE vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X656 a_3689_1685# a_3523_1685# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X662 temp1.dac.parallel_cells\[1\].vdac_batch.einvp_batch\[0\].pupd.TE a_5271_13647# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X669 vccd1 temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[3\].vref.TE a_4535_15823# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X684 vccd1 a_2623_1653# a_2539_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X690 a_7428_17607# temp1.capload\[5\].cap.TE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
R4 temp1.capload\[7\].cap_16.HI vccd1 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X691 a_2228_15095# a_2041_14735# a_2141_14851# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.107825 ps=1.36 w=0.42 l=0.15
X709 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref.TE _090_.A1 a_4418_16367# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X710 a_6600_15431# temp1.capload\[0\].cap_9.LO vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.32075 ps=1.685 w=0.42 l=0.15
X711 vccd1 _075_.A2 a_2877_14455# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.074375 ps=0.815 w=0.42 l=0.15
X712 vccd1 a_1766_2223# clkbuf_1_1__f_io_in[0].A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.14 ps=1.28 w=1 l=0.15
X720 vccd1 _065_.A a_2971_10383# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X724 vssd1 _093_.CLK a_1591_1685# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X730 vssd1 a_1674_2767# _093_.CLK vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X732 a_7084_15823# a_6835_15823# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X736 temp1.capload\[9\].cap.Z temp1.dcdc.Z a_7564_18319# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X741 a_2044_18319# temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref.TE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X742 vccd1 _051_.B1 a_4985_11177# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X747 a_7379_17705# temp1.dcdc.Z temp1.capload\[5\].cap.Z vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.27 ps=2.54 w=1 l=0.15
X750 vssd1 _095_.CLK a_3983_1135# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X752 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref.Z temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[4\].pupd.A a_1932_14441# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X753 vccd1 _048_.B a_2132_9295# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.3275 pd=1.655 as=0.195 ps=1.39 w=1 l=0.15
X755 vssd1 clkbuf_1_1__f_io_in[0].A a_1674_2767# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X762 vssd1 a_2932_21237# io_out[0] vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X763 vssd1 _075_.A2 a_3036_14197# vssd1 sky130_fd_pr__nfet_01v8 ad=0.122275 pd=1.08 as=0.05355 ps=0.675 w=0.42 l=0.15
X764 vssd1 a_4031_13866# input6.X vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X767 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref.Z temp1.dac.vdac_single.einvp_batch\[0\].pupd_20.HI a_20996_16143# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X770 vccd1 _048_.B a_3512_12559# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.3275 pd=1.655 as=0.195 ps=1.39 w=1 l=0.15
X777 a_2963_17231# temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref.Z temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref.Z vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.1755 ps=1.84 w=0.65 l=0.15
X778 temp1.capload\[6\].cap.Z temp1.dcdc.Z a_7084_15823# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X787 vssd1 del2.delay_chain\[3\].inv2.A a_3028_22691# vssd1 sky130_fd_pr__nfet_01v8 ad=0.14575 pd=1.63 as=0.05775 ps=0.76 w=0.55 l=0.15
X788 vssd1 temp1.dac.vdac_single.einvp_batch\[0\].vref_19.LO a_9135_16367# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X791 vccd1 a_2593_16413# a_2693_16631# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1085 ps=1.36 w=0.42 l=0.15
X794 vccd1 a_2927_11092# _057_.A1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X798 vssd1 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[4\].pupd.TE a_3063_18543# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X802 vccd1 temp1.dac.vdac_single.einvp_batch\[0\].pupd.TE a_20819_15823# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X810 vccd1 input6.X a_2406_12265# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1525 ps=1.305 w=1 l=0.15
X824 vccd1 a_1919_22325# _067_.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.26 ps=2.52 w=1 l=0.15
X826 a_5724_15279# temp1.dac.parallel_cells\[1\].vdac_batch.einvp_batch\[0\].pupd.TE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X832 vccd1 _111_.A _046_.B vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X833 _048_.B _111_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1425 ps=1.285 w=1 l=0.15
X836 a_8348_18231# temp1.capload\[1\].cap_10.LO vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.32075 ps=1.685 w=0.42 l=0.15
X839 io_out[1] a_1644_21781# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X846 a_2104_26677# _114_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X847 vssd1 a_5323_17973# temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[4\].pupd.TE vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.0567 ps=0.69 w=0.42 l=0.15
X857 a_1674_2767# clkbuf_1_1__f_io_in[0].A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=0.15
X866 a_4988_14441# _110_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.14825 ps=1.34 w=0.42 l=0.15
X868 vccd1 _069_.A a_2879_9839# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X875 a_4973_1135# a_3983_1135# a_4847_1501# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X877 vccd1 del2.delay_chain\[3\].inv2.A _046_.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.25
X885 vccd1 a_2455_3677# a_2623_3579# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X886 vccd1 _048_.A a_3983_20969# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X891 vssd1 _110_.A a_5271_14743# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X900 _095_.CLK a_1674_1135# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X903 a_2132_9295# _066_.A_N a_2041_9295# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.1525 ps=1.305 w=1 l=0.15
X908 a_2870_22691# del2.delay_chain\[3\].inv2.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.05775 pd=0.76 as=0.14575 ps=1.63 w=0.55 l=0.15
X909 vssd1 a_2238_13763# _090_.A2 vssd1 sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.08775 ps=0.92 w=0.65 l=0.15
X910 a_2229_9839# a_1959_10205# a_2139_10205# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X916 a_3791_17231# temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref.Z temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref.Z vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.1755 ps=1.84 w=0.65 l=0.15
X917 a_4712_16143# temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[3\].vref.TE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X918 a_4307_12167# a_4579_11995# a_4537_12265# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X923 a_2594_19631# del1.delay_chain\[3\].inv2.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.05775 pd=0.76 as=0.14575 ps=1.63 w=0.55 l=0.15
X924 vccd1 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref.TE a_1867_17455# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
R5 temp1.dac.vdac_single.einvp_batch\[0\].vref_19.LO vssd1 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X927 vssd1 a_2927_11092# _057_.A1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X935 vssd1 a_1674_1135# _095_.CLK vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X939 vssd1 temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[1\].pupd.TE a_4535_17455# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X940 vssd1 _060_.B a_4627_14191# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
X945 _072_.C_N a_2132_9295# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X950 vccd1 _115_.A _051_.A2 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X952 a_4590_1247# a_4422_1501# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X956 vccd1 io_in[1] a_1591_3855# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X957 vccd1 _051_.A2 a_3615_21263# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1475 pd=1.295 as=0.265 ps=2.53 w=1 l=0.15
X965 _046_.A del2.delay_chain\[3\].inv2.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.25
X966 a_4159_19087# _051_.Y temp1.dcdc.Z vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.27 ps=2.54 w=1 l=0.15
X967 a_4618_15055# _080_.A2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.095875 pd=0.945 as=0.17225 ps=1.83 w=0.65 l=0.15
X971 clkbuf_1_1__f_io_in[0].A a_1766_2223# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X977 a_3065_12021# _072_.C_N vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X989 _093_.CLK a_1674_2767# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X992 a_2104_25045# _113_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X996 vssd1 temp1.dcdc.Z temp1.inv2.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X997 a_1715_8779# _048_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X1001 a_4776_14165# a_4627_14191# a_5072_14441# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1006 a_2139_10205# a_1959_10205# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X1008 vccd1 temp1.capload\[7\].cap.TE a_6559_14735# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X1009 a_2030_3677# a_1757_3311# a_1945_3311# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X1012 _048_.B a_3983_18543# a_4171_18543# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1013 _085_.A1 a_4263_13109# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0.10025 ps=0.985 w=0.65 l=0.15
X1034 vssd1 del1.delay_chain\[2\].inv2.A del1.delay_chain\[2\].inv2.Y vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1040 clkbuf_1_1__f_io_in[0].A a_1766_2223# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X1046 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref.Z temp1.dac.parallel_cells\[1\].vdac_batch.einvp_batch\[0\].pupd.A a_5724_15279# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X1052 a_2104_25045# _113_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X1061 vssd1 a_1766_2223# clkbuf_1_1__f_io_in[0].A vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1071 a_4985_11177# _072_.C_N temp1.dac.parallel_cells\[0\].vdac_batch.einvp_batch\[0\].pupd.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X1073 _109_.A a_3983_10927# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1074 _093_.CLK a_1674_2767# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1077 a_2481_21807# _048_.A a_2409_21807# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X1078 temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[3\].vref.TE _085_.A1 a_4530_15279# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.089375 ps=0.925 w=0.65 l=0.15
X1080 _046_.A del2.delay_chain\[3\].inv2.A a_2870_22691# vssd1 sky130_fd_pr__nfet_01v8 ad=0.077 pd=0.83 as=0.05775 ps=0.76 w=0.55 l=0.15
X1085 del2.delay_chain\[0\].inv2.A del2.delay_chain\[0\].inv1.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1094 vccd1 a_2198_3423# a_2125_3677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X1098 vssd1 _109_.A temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref.TE vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X1101 _095_.CLK a_1674_1135# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1102 _048_.A del1.delay_chain\[3\].inv2.A a_2594_19631# vssd1 sky130_fd_pr__nfet_01v8 ad=0.077 pd=0.83 as=0.05775 ps=0.76 w=0.55 l=0.15
X1104 vccd1 _091_.A_N a_3983_10927# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X1108 a_3971_1679# a_3689_1685# a_3877_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0672 ps=0.74 w=0.42 l=0.15
X1113 vccd1 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[4\].pupd.TE a_1683_14191# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X1114 temp1.dac.parallel_cells\[0\].vdac_batch.einvp_batch\[0\].vref.TE _075_.A1 a_5722_14191# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.095875 ps=0.945 w=0.65 l=0.15
X1121 vssd1 a_3983_10927# _109_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X1123 _075_.A2 a_3065_12021# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.101875 ps=0.99 w=0.65 l=0.15
X1124 vssd1 temp1.capload\[3\].cap_12.LO a_7011_16367# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.235625 ps=1.375 w=0.65 l=0.15
X1125 a_2137_12879# _048_.B a_1919_12791# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X1127 vccd1 a_2840_26677# io_out[6] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X1136 vccd1 temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[3\].vref.TE a_5547_16367# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X1142 a_2840_26677# _115_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X1149 a_2125_3677# a_1591_3311# a_2030_3677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X1151 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref.Z temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref.Z a_4712_16143# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X1152 _090_.A2 a_2238_13763# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.101875 ps=0.99 w=0.65 l=0.15
X1154 vssd1 temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[3\].vref.TE a_3791_17231# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.235625 ps=1.375 w=0.65 l=0.15
X1157 a_7656_14191# temp1.dac.parallel_cells\[0\].vdac_batch.einvp_batch\[0\].vref.TE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X1165 a_4443_15529# _085_.A2 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1166 a_2321_10703# _048_.B a_2103_10615# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X1175 a_5796_17705# a_5547_17455# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X1179 vssd1 _079_.B a_4579_11995# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X1182 a_2927_9514# io_in[4] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X1185 _051_.Y _046_.B a_3698_21583# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.095875 ps=0.945 w=0.65 l=0.15
X1186 a_5447_18543# temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[1\].pupd.A temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref.Z vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.1755 ps=1.84 w=0.65 l=0.15
X1188 vssd1 _076_.X a_6559_13647# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X1190 a_2723_11791# _109_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X1200 vccd1 _075_.A2 a_5639_14441# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1475 pd=1.295 as=0.265 ps=2.53 w=1 l=0.15
X1208 vssd1 clkbuf_1_1__f_io_in[0].A a_1674_2767# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1209 a_1932_14441# a_1683_14191# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X1211 a_2139_10927# _111_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1013 ps=0.99 w=0.42 l=0.15
X1219 a_5496_18695# temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[1\].pupd.TE vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.32075 ps=1.685 w=0.42 l=0.15
X1220 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref.Z temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref.Z a_5796_17705# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X1225 vccd1 a_2011_10901# _063_.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.26 ps=2.52 w=1 l=0.15
X1226 vssd1 _079_.C a_3065_12021# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1230 vssd1 _066_.A_N a_2321_12015# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10075 ps=0.96 w=0.65 l=0.15
X1251 vssd1 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[4\].pupd.TE a_1591_13103# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X1265 vssd1 _111_.A a_2481_21807# vssd1 sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X1267 a_3983_20969# _048_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1278 vccd1 a_5271_14743# _051_.B1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X1279 vssd1 temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[1\].pupd.TE a_4619_17231# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.235625 ps=1.375 w=0.65 l=0.15
X1292 vccd1 temp1.dac.parallel_cells\[1\].vdac_batch.einvp_batch\[0\].pupd.TE a_5547_15823# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X1295 vssd1 a_1828_23957# io_out[3] vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X1298 _095_.CLK a_1674_1135# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1302 a_4668_17143# temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[1\].pupd.TE vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.32075 ps=1.685 w=0.42 l=0.15
X1303 vssd1 temp1.capload\[6\].cap_15.LO a_6835_15823# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X1304 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref.Z temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[4\].pupd.A a_2944_15529# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X1308 _109_.A a_3983_10927# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.07035 ps=0.755 w=0.42 l=0.15
X1309 vccd1 temp1.inv2.A _066_.B vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1322 vssd1 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[4\].pupd.TE a_3063_15823# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X1324 vssd1 del1.delay_chain\[3\].inv2.A a_2752_19631# vssd1 sky130_fd_pr__nfet_01v8 ad=0.14575 pd=1.63 as=0.05775 ps=0.76 w=0.55 l=0.15
X1326 vccd1 _046_.A a_3983_20969# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.385 ps=1.77 w=1 l=0.15
X1327 a_3331_19407# temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[4\].pupd.A temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref.Z vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.1755 ps=1.84 w=0.65 l=0.15
X1332 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref.Z temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[4\].pupd.A a_3240_18543# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X1335 vssd1 a_1766_2223# clkbuf_1_1__f_io_in[0].A vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1338 a_3893_14735# _051_.B1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1341 _109_.A a_3983_10927# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1342 vccd1 temp1.capload\[9\].cap.TE a_7387_17999# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X1345 a_3240_17455# temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[4\].pupd.TE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X1346 vccd1 a_2104_25045# io_out[4] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X1353 a_1945_1679# _063_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X1360 vssd1 a_2623_1653# a_2581_2057# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1368 _095_.CLK a_1674_1135# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1369 _091_.A_N a_2623_3579# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1384 a_2044_17455# temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref.TE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X1387 del2.delay_chain\[1\].inv2.Y del2.delay_chain\[1\].inv2.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1388 a_2576_19087# a_2327_19087# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X1389 vssd1 del2.delay_chain\[1\].inv1.A del2.delay_chain\[1\].inv2.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1392 vccd1 a_2007_11690# _063_.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X1394 vssd1 a_1674_1135# _095_.CLK vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1395 vccd1 a_3983_10927# _109_.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X1397 vssd1 a_1736_23413# io_out[2] vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X1399 vssd1 a_5015_1403# a_4973_1135# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1409 a_1757_1685# a_1591_1685# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1411 a_7011_16367# temp1.dcdc.Z temp1.capload\[3\].cap.Z vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.1755 ps=1.84 w=0.65 l=0.15
X1413 vccd1 a_1766_2223# clkbuf_1_1__f_io_in[0].A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1414 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref.TE _109_.A a_3984_16617# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1415 a_3204_13879# _110_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.101875 ps=0.99 w=0.42 l=0.15
X1419 vssd1 a_1674_2767# _093_.CLK vssd1 sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X1424 _069_.A a_1715_8779# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.16655 ps=1.39 w=1 l=0.15
X1431 temp1.dac.parallel_cells\[0\].vdac_batch.einvp_batch\[0\].vref.TE _109_.A a_5639_14441# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X1433 clkbuf_1_1__f_io_in[0].A a_1766_2223# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1434 vssd1 _115_.A a_2723_11791# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X1446 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref.Z temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref.Z a_2576_19087# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X1451 a_6551_15529# temp1.dcdc.Z temp1.capload\[0\].cap.Z vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.27 ps=2.54 w=1 l=0.15
X1459 _085_.A2 a_2421_13109# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.14825 ps=1.34 w=1 l=0.15
X1464 a_3984_16617# _109_.A temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref.TE vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.14 ps=1.28 w=1 l=0.15
X1467 vccd1 a_2104_26677# io_out[5] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X1468 vssd1 del1.delay_chain\[2\].inv1.A del1.delay_chain\[2\].inv2.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1469 a_4345_13353# a_4157_13149# a_4263_13109# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X1473 a_6784_17143# temp1.capload\[8\].cap.TE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X1475 _087_.A a_2233_15939# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X1481 _046_.B _048_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1490 a_3012_17143# temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[3\].vref.TE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X1491 a_2406_12265# _066_.A_N a_2103_11989# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1525 pd=1.305 as=0.195 ps=1.39 w=1 l=0.15
X1492 _093_.CLK a_1674_2767# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1496 vccd1 a_3983_18543# _048_.B vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1497 a_7428_18695# temp1.capload\[4\].cap_13.LO vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.32075 ps=1.685 w=0.42 l=0.15
X1498 vccd1 a_1674_1135# _095_.CLK vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.14 ps=1.28 w=1 l=0.15
X1499 _053_.A1 a_1591_7663# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X1501 vccd1 del2.delay_chain\[3\].inv2.A _046_.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.25
X1503 vssd1 _110_.A a_2238_13763# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X1508 vssd1 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref.TE a_2327_19087# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X1509 _048_.B _111_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1510 temp1.dac.vdac_single.einvp_batch\[0\].pupd.TE _071_.C a_3977_14735# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
R6 vccd1 temp1.dac.vdac_single.einvp_batch\[0\].vref_19.HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X1520 vccd1 a_6600_15431# a_6551_15529# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1825 ps=1.365 w=1 l=0.15
X1525 a_4208_19319# temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref.Z vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.32075 ps=1.685 w=0.42 l=0.15
X1536 _051_.B1 a_5271_14743# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X1540 vssd1 _083_.C_N temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[1\].pupd.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1543 _065_.A a_2139_10205# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X1547 a_5724_16143# temp1.dac.parallel_cells\[1\].vdac_batch.einvp_batch\[0\].pupd.TE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X1549 vccd1 a_4307_12167# _080_.A1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.275 ps=2.55 w=1 l=0.15
X1554 io_out[3] a_1828_23957# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X1557 a_1959_9615# _066_.A_N vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.08775 ps=0.92 w=0.65 l=0.15
X1562 a_2927_9514# io_in[4] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1564 vssd1 io_in[1] a_1591_3855# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X1568 a_7428_17607# temp1.capload\[5\].cap.TE vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.32075 ps=1.685 w=0.42 l=0.15
X1569 temp1.capload\[7\].cap.Z temp1.dcdc.Z a_6808_14735# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X1573 vccd1 a_4558_1653# _111_.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1425 pd=1.285 as=0.135 ps=1.27 w=1 l=0.15
X1580 vssd1 temp1.dac.parallel_cells\[1\].vdac_batch.einvp_batch\[1\].vref.TE a_5547_17455# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X1582 a_3345_13353# _051_.B1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X1587 a_3219_12265# _072_.C_N a_3147_12265# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X1590 a_2133_15823# _109_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.10785 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X1597 a_2198_1653# a_2030_1679# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X1600 _109_.A a_3983_10927# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X1604 a_2593_23145# _048_.B _112_.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X1605 _111_.A a_4558_1653# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.105625 ps=0.975 w=0.65 l=0.15
X1609 _051_.A2 _048_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1610 vccd1 a_1674_2767# _093_.CLK vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.14 ps=1.28 w=1 l=0.15
X1614 vssd1 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[4\].pupd.TE a_1683_14191# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X1626 a_3840_17143# temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[3\].vref.TE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X1637 vccd1 _085_.A2 a_4443_15529# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.28 ps=2.56 w=1 l=0.15
X1639 io_out[2] a_1736_23413# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X1641 vssd1 _051_.B1 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[4\].pupd.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X1643 a_1644_21781# _110_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X1650 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref.TE _109_.A a_3984_16617# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.26 ps=2.52 w=1 l=0.15
X1655 temp1.dac.parallel_cells\[1\].vdac_batch.einvp_batch\[1\].vref.TE _109_.A a_4535_14735# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X1660 vccd1 temp1.dac.vdac_single.einvp_batch\[0\].vref_19.LO a_9135_16367# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X1662 vccd1 a_2455_1679# a_2623_1653# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1665 clkbuf_1_1__f_io_in[0].A a_1766_2223# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1673 a_4471_1679# a_3689_1685# a_4387_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.09135 pd=0.855 as=0.0567 ps=0.69 w=0.42 l=0.15
X1687 vccd1 a_3204_13879# _080_.A2 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.28 ps=2.56 w=1 l=0.15
X1688 a_5353_12265# _079_.B temp1.dac.parallel_cells\[1\].vdac_batch.einvp_batch\[0\].pupd.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X1692 vssd1 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref.Z a_4159_19407# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.235625 ps=1.375 w=0.65 l=0.15
X1699 a_2693_16631# _090_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.074375 pd=0.815 as=0.0567 ps=0.69 w=0.42 l=0.15
X1700 a_2455_3677# a_1591_3311# a_2198_3423# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X1704 a_1766_2223# io_in[0] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1705 a_4517_1501# a_3983_1135# a_4422_1501# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X1706 vssd1 a_4847_1501# a_5015_1403# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1711 a_5496_18695# temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[1\].pupd.TE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X1713 a_1736_23413# _111_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X1717 a_3983_20969# _115_.A _066_.A_N vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1723 vccd1 a_2103_10615# _079_.B vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.3275 pd=1.655 as=0.28 ps=2.56 w=1 l=0.15
X1726 vccd1 _111_.A _048_.B vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1727 a_2777_14237# _109_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1087 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X1733 vccd1 a_2095_22657# a_1919_22325# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.0609 ps=0.71 w=0.42 l=0.15
X1734 vccd1 a_1644_21781# io_out[1] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X1735 vccd1 a_1674_1135# _095_.CLK vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1745 del2.delay_chain\[2\].inv2.Y del2.delay_chain\[2\].inv2.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1748 vccd1 _048_.A a_3983_20969# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.145 ps=1.29 w=1 l=0.15
X1750 _095_.CLK a_1674_1135# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1754 a_2828_20407# temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref.TE vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.32075 ps=1.685 w=0.42 l=0.15
X1756 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref.Z temp1.dac.parallel_cells\[1\].vdac_batch.einvp_batch\[0\].pupd.A a_5724_16143# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X1761 vccd1 _048_.A a_2593_23145# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X1762 a_2944_15529# a_2695_15279# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
R7 vssd1 temp1.capload\[0\].cap_9.LO sky130_fd_pr__res_generic_po w=0.48 l=0.045
X1777 a_1920_28853# _116_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X1780 vccd1 _081_.X a_5271_13647# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X1782 _068_.B a_1591_6031# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X1784 a_6735_17231# temp1.dcdc.Z temp1.capload\[8\].cap.Z vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.1755 ps=1.84 w=0.65 l=0.15
X1787 vssd1 a_2103_11989# _060_.B vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1789 vccd1 temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[1\].pupd.TE a_4535_17455# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X1791 a_2041_9295# _053_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1525 pd=1.305 as=0.26 ps=2.52 w=1 l=0.15
X1796 a_1919_22325# a_2095_22657# a_2047_22717# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0504 ps=0.66 w=0.42 l=0.15
X1798 vccd1 a_2623_3579# a_2539_3677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X1802 a_4443_15529# _109_.A temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[3\].vref.TE vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.36 pd=2.72 as=0.135 ps=1.27 w=1 l=0.15
X1803 a_2198_3423# a_2030_3677# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X1804 a_4418_16367# _090_.A2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X1812 _095_.CLK a_1674_1135# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X1818 a_3512_12559# _048_.B a_3339_12879# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X1827 _053_.A1 a_1591_7663# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1832 vccd1 a_1674_2767# _093_.CLK vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1837 vssd1 a_1674_1135# _095_.CLK vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1838 vccd1 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[4\].pupd.TE a_1591_13103# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X1841 a_7980_13879# temp1.dac.parallel_cells\[0\].vdac_batch.einvp_batch\[0\].pupd.TE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X1845 a_2137_12879# _057_.A1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1849 a_2198_1653# a_2030_1679# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X1851 vssd1 _090_.A2 a_4418_16367# vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X1853 a_3036_14197# _075_.A1 a_2964_14197# vssd1 sky130_fd_pr__nfet_01v8 ad=0.05355 pd=0.675 as=0.0441 ps=0.63 w=0.42 l=0.15
R8 temp1.capload\[6\].cap_15.HI vccd1 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X1857 vssd1 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[4\].pupd.TE a_3155_17999# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X1866 clkbuf_1_1__f_io_in[0].A a_1766_2223# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1867 a_2455_1679# a_1757_1685# a_2198_1653# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1869 del1.delay_chain\[1\].inv1.Y del1.delay_chain\[1\].inv1.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1872 a_2503_13353# _079_.C a_2421_13109# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X1876 a_1945_3311# _061_.B1_N vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X1878 del1.delay_chain\[3\].inv2.A del1.delay_chain\[2\].inv2.Y vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1879 _068_.B a_1591_6031# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1882 _048_.B a_3983_18543# a_4171_18543# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1897 clkbuf_1_1__f_io_in[0].A a_1766_2223# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1902 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref.Z temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[4\].pupd.A a_3332_18319# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X1903 vccd1 a_3012_17143# a_2963_16911# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1825 ps=1.365 w=1 l=0.15
X1905 a_4171_18543# a_3983_18543# _048_.B vssd1 sky130_fd_pr__nfet_01v8 ad=0.092625 pd=0.935 as=0.08775 ps=0.92 w=0.65 l=0.15
X1906 a_7728_14441# a_7479_14191# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X1907 io_out[1] a_1644_21781# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X1908 a_3983_20969# _111_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1913 _093_.CLK a_1674_2767# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X1915 vccd1 _093_.CLK a_1591_3311# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1922 vccd1 _051_.B1 a_4417_13353# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.06825 ps=0.745 w=0.42 l=0.15
X1926 vccd1 _090_.A2 a_2693_16631# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.074375 ps=0.815 w=0.42 l=0.15
X1930 a_1840_13353# a_1591_13103# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X1934 _066_.A_N _115_.A a_3983_20969# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.32 ps=2.64 w=1 l=0.15
X1938 vccd1 a_4776_14165# _090_.A1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.135 ps=1.27 w=1 l=0.15
X1947 vccd1 a_2133_15823# a_2233_15939# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1085 ps=1.36 w=0.42 l=0.15
X1955 a_7428_18695# temp1.capload\[4\].cap_13.LO vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X1958 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref.Z temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref.Z a_1932_16617# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X1960 vssd1 a_4558_1653# _111_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.08775 ps=0.92 w=0.65 l=0.15
X1963 a_3983_20969# _115_.A _066_.A_N vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.385 pd=1.77 as=0.135 ps=1.27 w=1 l=0.15
X1973 vccd1 _046_.A a_3983_20969# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1977 io_out[4] a_2104_25045# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X1982 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref.Z temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[4\].pupd.A a_1840_13353# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X1992 vssd1 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref.TE a_2779_20495# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.235625 ps=1.375 w=0.65 l=0.15
X1995 vssd1 a_4558_1653# a_4516_2057# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1197 pd=1.41 as=0.066 ps=0.745 w=0.42 l=0.15
X1997 vssd1 a_1766_2223# clkbuf_1_1__f_io_in[0].A vssd1 sky130_fd_pr__nfet_01v8 ad=0.05775 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X2005 vssd1 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref.TE a_1867_15279# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X2015 a_2409_21807# _046_.A a_2327_21807# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X2016 vccd1 a_7428_18695# a_7379_18793# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1825 ps=1.365 w=1 l=0.15
X2019 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref.Z temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref.Z a_2044_15279# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X2020 vccd1 _110_.A a_3219_12265# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X2028 vccd1 del1.delay_chain\[0\].inv2.A del1.delay_chain\[1\].inv1.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X2032 vssd1 a_2455_1679# a_2623_1653# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2034 a_4418_16367# _090_.A1 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref.TE vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X2037 temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[3\].vref.TE _109_.A a_4443_15529# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2041 vssd1 _051_.B1 a_4263_13109# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X2042 a_2116_17999# a_1867_17999# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X2043 a_2575_13353# _083_.C_N a_2503_13353# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X2049 a_2539_1679# a_1757_1685# a_2455_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X2050 vssd1 a_1674_2767# _093_.CLK vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2073 a_4149_1135# a_3983_1135# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2075 io_out[5] a_2104_26677# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X2078 vccd1 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref.TE a_1867_17999# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X2079 vssd1 _066_.A_N a_2137_12879# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10075 ps=0.96 w=0.65 l=0.15
X2091 a_5724_16367# temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[3\].vref.TE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X2092 temp1.dac.parallel_cells\[1\].vdac_batch.einvp_batch\[0\].pupd.TE a_5271_13647# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2093 vccd1 _061_.B1_N a_1959_10205# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X2098 a_4350_11587# _051_.B1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.14825 ps=1.34 w=0.42 l=0.15
X2099 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref.Z temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref.Z a_2116_17999# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X2101 a_4590_1247# a_4422_1501# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X2104 a_3877_1679# _065_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.1092 ps=1.36 w=0.42 l=0.15
X2106 a_3312_17705# a_3063_17455# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X2108 a_2320_13763# _079_.C a_2238_13763# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X2110 a_2321_12015# input6.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2112 vccd1 _046_.A a_3983_18543# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X2123 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[4\].pupd.TE a_5323_17973# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2133 vssd1 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref.TE a_3607_20495# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.235625 ps=1.375 w=0.65 l=0.15
X2134 vssd1 _111_.A a_4171_18543# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.092625 ps=0.935 w=0.65 l=0.15
X2135 a_2327_21807# _048_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X2136 a_2030_1679# a_1591_1685# a_1945_1679# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
R9 vssd1 temp1.capload\[1\].cap_10.LO sky130_fd_pr__res_generic_po w=0.48 l=0.045
X2142 vssd1 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[4\].pupd.TE a_2695_15279# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X2146 input7.X a_1591_13647# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X2147 temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[1\].pupd.A _051_.B1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2151 a_2116_17705# a_1867_17455# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X2153 a_1766_2223# io_in[0] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X2159 vccd1 _111_.A a_3983_20969# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2160 temp1.dac.parallel_cells\[0\].vdac_batch.einvp_batch\[0\].pupd.A _072_.C_N vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2162 a_4576_18231# temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[1\].pupd.TE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X2168 del1.delay_chain\[2\].inv1.A del1.delay_chain\[1\].inv1.Y vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X2170 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref.Z temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[4\].pupd.A a_3312_17705# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X2176 a_4619_17231# temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[1\].pupd.A temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref.Z vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.1755 ps=1.84 w=0.65 l=0.15
X2179 vssd1 _091_.A_N a_3983_10927# vssd1 sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.1113 ps=1.37 w=0.42 l=0.15
X2181 a_20996_16143# temp1.dac.vdac_single.einvp_batch\[0\].pupd.TE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X2182 vccd1 a_1674_1135# _095_.CLK vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2183 vccd1 _072_.C_N a_4487_11561# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X2185 a_4413_20719# _048_.A a_4771_20719# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2188 io_out[0] a_2932_21237# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X2190 _090_.A1 a_4776_14165# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14575 ps=1.335 w=1 l=0.15
X2191 _081_.X a_2141_14851# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X2192 a_2964_14197# a_2777_14237# a_2877_14455# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.107825 ps=1.36 w=0.42 l=0.15
X2198 a_2156_2057# a_1757_1685# a_2030_1679# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X2199 _095_.CLK a_1674_1135# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2202 a_7931_13967# temp1.dac.parallel_cells\[0\].vdac_batch.einvp_batch\[0\].pupd.A temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref.Z vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.1755 ps=1.84 w=0.65 l=0.15
X2203 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref.Z temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref.Z a_2116_17705# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X2205 vccd1 a_8348_18231# a_8299_17999# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1825 ps=1.365 w=1 l=0.15
R10 temp1.capload\[5\].cap_14.HI vccd1 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X2207 vccd1 temp1.dac.parallel_cells\[0\].vdac_batch.einvp_batch\[0\].vref.TE a_7479_14191# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X2213 a_3983_20969# _046_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2217 a_1757_1685# a_1591_1685# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2221 _093_.CLK a_1674_2767# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2226 a_3977_14735# _109_.A a_3893_14735# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2234 vssd1 temp1.capload\[5\].cap.TE a_7379_17455# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.235625 ps=1.375 w=0.65 l=0.15
X2242 a_2517_23439# _046_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X2247 a_4149_1135# a_3983_1135# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2249 a_4847_1501# a_3983_1135# a_4590_1247# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X2253 _051_.A2 _115_.A a_3333_20719# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2254 a_3028_22691# del2.delay_chain\[3\].inv2.A _046_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.05775 pd=0.76 as=0.077 ps=0.83 w=0.55 l=0.15
X2259 a_4537_12265# _071_.C a_4442_12265# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.06825 ps=0.745 w=0.42 l=0.15
X2271 _092_.A a_2693_16631# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.122275 ps=1.08 w=0.65 l=0.15
X2273 a_4418_16367# _090_.A1 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref.TE vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X2274 _111_.A a_4558_1653# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1425 ps=1.285 w=1 l=0.15
X2275 a_4527_17999# temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[1\].pupd.A temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref.Z vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.27 ps=2.54 w=1 l=0.15
X2276 vccd1 del2.delay_chain\[0\].inv2.A del2.delay_chain\[1\].inv1.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X2278 vccd1 a_1674_2767# _093_.CLK vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2283 a_2392_13763# _060_.B a_2320_13763# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X2284 a_4263_13109# _071_.C vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X2286 a_2041_14735# _109_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.10785 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X2288 vssd1 a_2011_10901# _063_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.169 ps=1.82 w=0.65 l=0.15
X2314 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref.Z temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref.Z a_5724_16367# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X2321 a_3380_19319# temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[4\].pupd.TE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X2328 a_2593_16413# _091_.A_N vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.10785 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X2334 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref.Z temp1.dac.vdac_single.einvp_batch\[0\].pupd_20.HI a_21068_15823# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X2337 clkbuf_1_1__f_io_in[0].A a_1766_2223# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.05775 ps=0.695 w=0.42 l=0.15
X2338 a_3984_16617# _090_.A2 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2342 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref.Z temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref.Z a_7728_14441# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X2343 a_2963_16911# temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref.Z temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref.Z vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.27 ps=2.54 w=1 l=0.15
R11 vssd1 temp1.dac.vdac_single.einvp_batch\[0\].pupd_20.LO sky130_fd_pr__res_generic_po w=0.48 l=0.045
X2348 _091_.A_N a_2623_3579# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2352 vccd1 _046_.A a_2327_21807# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2354 vccd1 _111_.A _048_.B vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.39 pd=2.78 as=0.135 ps=1.27 w=1 l=0.15
X2361 vssd1 temp1.capload\[2\].cap.TE a_7755_16367# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X2368 vssd1 temp1.inv2.A _066_.B vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2369 a_6736_15055# temp1.capload\[7\].cap.TE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X2371 a_3656_20407# temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref.TE vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.32075 ps=1.685 w=0.42 l=0.15
X2376 a_2103_10615# _048_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.3275 ps=1.655 w=1 l=0.15
X2378 temp1.capload\[2\].cap.Z temp1.dcdc.Z a_7932_16367# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X2384 vccd1 temp1.dac.parallel_cells\[1\].vdac_batch.einvp_batch\[1\].vref.TE a_5547_17455# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X2388 a_4215_11703# a_4487_11561# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2400 _093_.CLK a_1674_2767# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2402 _113_.A _046_.B a_2517_23439# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X2405 a_1932_16617# a_1683_16367# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X2408 vccd1 a_4215_11703# _075_.A1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.275 ps=2.55 w=1 l=0.15
X2411 _079_.C _048_.B a_4259_12879# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2422 _095_.CLK a_1674_1135# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2439 del2.delay_chain\[1\].inv2.Y del2.delay_chain\[1\].inv2.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2445 a_1674_1135# clkbuf_1_1__f_io_in[0].A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2450 vccd1 _080_.A2 a_2141_14851# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.074375 ps=0.815 w=0.42 l=0.15
X2452 vccd1 a_1766_2223# clkbuf_1_1__f_io_in[0].A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2453 a_1945_3311# _061_.B1_N vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X2455 a_2877_14455# _075_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.074375 pd=0.815 as=0.0567 ps=0.69 w=0.42 l=0.15
X2456 vssd1 a_5015_1403# _110_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2464 a_3791_16911# temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref.Z temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref.Z vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.27 ps=2.54 w=1 l=0.15
X2469 vccd1 a_2187_10901# a_2011_10901# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.0609 ps=0.71 w=0.42 l=0.15
X2470 vssd1 _060_.B temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[4\].pupd.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2473 vccd1 _068_.B a_1715_8779# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
R12 vccd1 temp1.capload\[9\].cap_18.HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X2475 vccd1 io_in[0] a_1766_2223# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2478 vssd1 a_1674_2767# _093_.CLK vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2488 a_6239_18708# _087_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X2491 vssd1 temp1.capload\[0\].cap_9.LO a_6551_15279# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.235625 ps=1.375 w=0.65 l=0.15
X2493 _076_.X a_2877_14455# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X2502 vccd1 _110_.A a_2575_13353# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X2504 vssd1 _051_.B1 temp1.dac.parallel_cells\[0\].vdac_batch.einvp_batch\[0\].pupd.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2510 vccd1 a_3840_17143# a_3791_16911# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1825 ps=1.365 w=1 l=0.15
X2514 vccd1 _080_.A2 a_4535_14735# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1475 pd=1.295 as=0.265 ps=2.53 w=1 l=0.15
X2516 _093_.CLK a_1674_2767# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2521 vccd1 temp1.dac.parallel_cells\[1\].vdac_batch.einvp_batch\[1\].vref.TE a_5547_16911# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X2525 _116_.A a_1959_27247# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X2526 a_4771_20719# _048_.A a_4413_20719# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2528 vccd1 a_2932_21237# io_out[0] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X2530 a_3983_20969# _111_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
R13 vccd1 temp1.capload\[2\].cap_11.HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X2533 a_1674_2767# clkbuf_1_1__f_io_in[0].A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2539 vssd1 a_4387_1679# a_4558_1653# vssd1 sky130_fd_pr__nfet_01v8 ad=0.105625 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X2540 a_4159_19407# _051_.Y temp1.dcdc.Z vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.1755 ps=1.84 w=0.65 l=0.15
X2544 vssd1 input7.X a_4259_12879# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X2547 a_3984_16617# _090_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2553 vccd1 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref.TE a_1591_16911# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X2558 _066_.A_N _115_.A a_3983_20969# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2564 a_9312_16367# temp1.dac.vdac_single.einvp_batch\[0\].vref_19.LO vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X2565 a_6808_14735# a_6559_14735# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X2567 vssd1 _061_.B1_N a_2187_10901# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X2568 a_3240_18543# temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[4\].pupd.TE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X2581 a_3983_20969# _048_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2595 a_4701_15279# _085_.A1 temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[3\].vref.TE vssd1 sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.091 ps=0.93 w=0.65 l=0.15
X2607 a_5323_17973# _092_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.06825 ps=0.745 w=0.42 l=0.15
X2608 a_2752_19631# del1.delay_chain\[3\].inv2.A _048_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.05775 pd=0.76 as=0.077 ps=0.83 w=0.55 l=0.15
X2609 a_4784_15823# a_4535_15823# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X2616 vssd1 _071_.C a_4776_14165# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X2619 vccd1 a_4668_17143# a_4619_16911# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1825 ps=1.365 w=1 l=0.15
X2622 _095_.CLK a_1674_1135# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2624 a_1801_8779# _048_.A a_1715_8779# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X2628 vccd1 a_2041_14735# a_2141_14851# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1085 ps=1.36 w=0.42 l=0.15
X2631 vssd1 temp1.dac.parallel_cells\[0\].vdac_batch.einvp_batch\[0\].vref.TE a_7479_14191# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X2638 a_4031_13866# io_in[6] vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X2640 vccd1 a_4847_1501# a_5015_1403# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X2643 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref.Z temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[4\].pupd.A a_3240_16143# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X2644 a_4422_1501# a_4149_1135# a_4337_1135# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X2649 vccd1 a_2238_13763# _090_.A2 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.315 pd=2.63 as=0.135 ps=1.27 w=1 l=0.15
X2650 vccd1 a_1766_2223# clkbuf_1_1__f_io_in[0].A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X2653 vssd1 a_1766_2223# clkbuf_1_1__f_io_in[0].A vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2658 temp1.dac.parallel_cells\[0\].vdac_batch.einvp_batch\[0\].pupd.TE a_6559_13647# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X2661 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref.Z temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref.Z a_4784_15823# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X2662 vccd1 a_4576_18231# a_4527_17999# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1825 ps=1.365 w=1 l=0.15
X2667 vssd1 del2.delay_chain\[1\].inv2.Y del2.delay_chain\[2\].inv2.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2673 vssd1 temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[3\].vref.TE a_4535_15823# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X2679 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[4\].pupd.A _060_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2688 vssd1 _051_.B1 _051_.Y vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X2691 _085_.A2 a_2421_13109# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.101875 ps=0.99 w=0.65 l=0.15
X2694 vccd1 a_2927_9514# _055_.A1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X2701 a_4712_17455# temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[1\].pupd.TE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X2708 vccd1 _061_.B1_N a_2956_11445# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.18575 pd=1.415 as=0.1176 ps=1.4 w=0.42 l=0.15
X2709 vccd1 _060_.B a_4627_14191# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.1092 ps=1.36 w=0.42 l=0.15
X2714 a_4171_18543# a_3983_18543# _048_.B vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2718 vssd1 a_1674_1135# _095_.CLK vssd1 sky130_fd_pr__nfet_01v8 ad=0.05775 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X2723 vssd1 _111_.A a_4171_18543# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2728 a_2890_11471# a_2956_11445# a_2723_11791# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10725 ps=0.98 w=0.65 l=0.15
X2736 a_5724_17231# temp1.dac.parallel_cells\[1\].vdac_batch.einvp_batch\[1\].vref.TE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
R14 vccd1 temp1.capload\[3\].cap_12.HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X2737 vccd1 a_1674_1135# _095_.CLK vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2739 vssd1 a_1644_21781# io_out[1] vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X2740 vccd1 _111_.A a_3983_20969# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2741 vssd1 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref.TE a_1683_16367# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X2749 vccd1 a_4590_1247# a_4517_1501# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X2753 a_3984_16617# _090_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.145 ps=1.29 w=1 l=0.15
X2755 a_2504_19407# temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref.TE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X2760 io_out[7] a_1920_28853# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X2762 vssd1 _085_.A2 a_4701_15279# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.06825 ps=0.86 w=0.65 l=0.15
X2764 vccd1 a_2623_1653# _115_.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2765 vccd1 clkbuf_1_1__f_io_in[0].A a_1674_1135# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2767 vssd1 a_4307_12167# _080_.A1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.17875 ps=1.85 w=0.65 l=0.15
X2775 vssd1 _071_.C a_4307_12167# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X2779 clkbuf_1_1__f_io_in[0].A a_1766_2223# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2780 vccd1 _095_.CLK a_3523_1685# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X2786 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref.Z temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref.Z a_9312_16367# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X2789 a_1919_22325# _066_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.2279 ps=1.74 w=0.42 l=0.15
X2791 a_2233_15939# _085_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.074375 pd=0.815 as=0.0567 ps=0.69 w=0.42 l=0.15
X2796 vssd1 a_4130_1653# a_4068_2057# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1493 pd=1.22 as=0.0687 ps=0.76 w=0.42 l=0.15
X2804 vccd1 _051_.B1 a_2139_10205# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X2806 vccd1 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref.TE a_1867_15279# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X2808 _093_.CLK a_1674_2767# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2810 a_3983_20969# _046_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.135 ps=1.27 w=1 l=0.15
X2811 vssd1 temp1.dac.vdac_single.einvp_batch\[0\].pupd.TE a_20819_15823# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X2815 a_6239_18708# _087_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2827 a_3333_20719# _048_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2842 a_2779_20495# temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref.Z temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref.Z vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.1755 ps=1.84 w=0.65 l=0.15
X2843 a_2455_3677# a_1757_3311# a_2198_3423# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2844 a_3147_12265# _079_.C a_3065_12021# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X2845 vccd1 a_1674_2767# _093_.CLK vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2853 _116_.A a_1959_27247# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2858 a_1674_1135# clkbuf_1_1__f_io_in[0].A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X2863 vccd1 _055_.A1 a_2406_10383# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1525 ps=1.305 w=1 l=0.15
R15 temp1.dac.vdac_single.einvp_batch\[0\].pupd_20.HI vccd1 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X2865 vssd1 a_4157_13149# a_4263_13109# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2869 vccd1 clkbuf_1_1__f_io_in[0].A a_1674_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2876 vccd1 a_4130_1653# a_4064_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.0693 ps=0.75 w=0.42 l=0.15
X2881 vssd1 input7.X a_3339_12879# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2884 _090_.A2 a_2238_13763# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14825 ps=1.34 w=1 l=0.15
X2890 a_7060_16519# temp1.capload\[3\].cap_12.LO vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X2892 vccd1 a_1919_12791# _083_.C_N vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.3275 pd=1.655 as=0.28 ps=2.56 w=1 l=0.15
X2897 a_3204_13879# _079_.C a_3435_13763# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X2900 vssd1 a_1674_2767# _093_.CLK vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2902 vccd1 del2.delay_chain\[1\].inv1.A del2.delay_chain\[1\].inv2.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X2913 vssd1 _072_.C_N a_4487_11561# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X2917 _071_.C a_3512_12559# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.3275 ps=1.655 w=1 l=0.15
X2921 temp1.dac.parallel_cells\[1\].vdac_batch.einvp_batch\[0\].pupd.A _079_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2923 a_3615_21263# _046_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1475 ps=1.295 w=1 l=0.15
X2927 a_4157_13149# _083_.C_N vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X2930 a_2890_11471# _109_.A a_2818_11471# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.105 ps=1.21 w=1 l=0.15
X2932 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref.Z temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[1\].pupd.A a_4712_17455# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X2936 vccd1 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[4\].pupd.TE a_2695_15279# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X2940 temp1.dac.parallel_cells\[1\].vdac_batch.einvp_batch\[1\].vref.TE _080_.A1 a_4618_15055# vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.095875 ps=0.945 w=0.65 l=0.15
X2941 a_1766_2223# io_in[0] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2950 _066_.A_N _115_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2958 vccd1 a_5323_17973# temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[4\].pupd.TE vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X2961 a_1674_2767# clkbuf_1_1__f_io_in[0].A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X2963 a_4171_18543# _111_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2965 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref.Z temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref.Z a_5724_17231# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X2969 vssd1 a_1674_1135# _095_.CLK vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2970 a_3607_20495# temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref.Z temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref.Z vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.1755 ps=1.84 w=0.65 l=0.15
X2973 a_4413_20719# _046_.A _066_.A_N vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2975 vssd1 _071_.C a_4215_11703# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X2980 _079_.C _066_.A_N a_4341_12559# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.39 as=0.105 ps=1.21 w=1 l=0.15
X2988 a_4413_20719# _048_.A a_4771_20719# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2991 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref.Z temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref.Z a_2504_19407# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X2995 a_4530_15279# _085_.A2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.18525 ps=1.87 w=0.65 l=0.15
X2998 vccd1 a_7060_16519# a_7011_16617# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1825 ps=1.365 w=1 l=0.15
X3003 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref.Z temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref.Z a_1768_17231# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X3024 del2.delay_chain\[3\].inv2.A del2.delay_chain\[2\].inv2.Y vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X3047 a_7379_18793# temp1.dcdc.Z temp1.capload\[4\].cap.Z vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.27 ps=2.54 w=1 l=0.15
X3053 a_5796_15529# a_5547_15279# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X3057 vccd1 _110_.A a_5271_14743# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X3058 vssd1 a_2927_9514# _055_.A1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X3059 _065_.X a_2971_10383# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X3064 _095_.CLK a_1674_1135# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.05775 ps=0.695 w=0.42 l=0.15
X3067 a_1919_12791# _048_.B vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.3275 ps=1.655 w=1 l=0.15
X3072 a_7379_17455# temp1.dcdc.Z temp1.capload\[5\].cap.Z vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.1755 ps=1.84 w=0.65 l=0.15
X3075 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref.Z temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[4\].pupd.A a_1860_14191# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X3079 a_2133_15823# _109_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1087 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X3082 _115_.A a_2623_1653# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3090 _095_.CLK a_1674_1135# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3093 io_out[6] a_2840_26677# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X3097 a_8348_18231# temp1.capload\[1\].cap_10.LO vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X3098 vccd1 a_1766_2223# clkbuf_1_1__f_io_in[0].A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3102 vssd1 a_1919_12791# _083_.C_N vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X3105 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref.Z temp1.dac.parallel_cells\[1\].vdac_batch.einvp_batch\[0\].pupd.A a_5796_15529# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X3107 a_2030_3677# a_1591_3311# a_1945_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X3121 vccd1 io_in[0] a_1766_2223# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3122 a_2539_3677# a_1757_3311# a_2455_3677# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X3125 vccd1 a_1736_23413# io_out[2] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X3126 a_4443_15529# _085_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3129 a_3332_18319# temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[4\].pupd.TE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X3130 a_4847_1501# a_4149_1135# a_4590_1247# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X3137 a_3984_16617# _109_.A temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref.TE vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3139 a_2987_14735# _051_.B1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X3142 vssd1 a_1920_28853# io_out[7] vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X3147 vssd1 temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[1\].pupd.TE a_4527_18319# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.235625 ps=1.375 w=0.65 l=0.15
X3149 a_4771_20719# _111_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3150 vssd1 _081_.X a_5271_13647# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X3152 vssd1 a_2623_1653# _115_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3158 a_5639_14441# _075_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1475 ps=1.295 w=1 l=0.15
X3159 a_2156_3311# a_1757_3311# a_2030_3677# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X3162 vccd1 a_2777_14237# a_2877_14455# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1085 ps=1.36 w=0.42 l=0.15
X3166 a_2321_12015# _048_.B a_2103_11989# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X3168 vccd1 temp1.capload\[2\].cap.TE a_7755_16367# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X3179 vssd1 _115_.A _066_.A_N vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.208 ps=1.94 w=0.65 l=0.15
X3180 vssd1 temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[1\].pupd.TE a_5447_18543# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.235625 ps=1.375 w=0.65 l=0.15
X3181 _093_.CLK a_1674_2767# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3184 vccd1 del1.delay_chain\[2\].inv1.A del1.delay_chain\[2\].inv2.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X3193 vccd1 io_in[7] a_1591_13647# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X3199 _066_.A_N _115_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3204 a_4215_11703# _051_.B1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.10025 ps=0.985 w=0.42 l=0.15
X3205 a_8299_17999# temp1.dcdc.Z temp1.capload\[1\].cap.Z vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.27 ps=2.54 w=1 l=0.15
X3207 vccd1 clkbuf_1_1__f_io_in[0].A a_1674_1135# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3208 vccd1 _111_.A a_2327_21807# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.142225 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X3209 a_5796_15823# a_5547_15823# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X3210 vssd1 a_2198_3423# a_2156_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X3219 vccd1 a_5496_18695# a_5447_18793# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1825 ps=1.365 w=1 l=0.15
X3227 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref.Z temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[4\].pupd.A a_1768_13103# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X3240 _093_.CLK a_1674_2767# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3241 a_4068_2057# a_3689_1685# a_3971_1679# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0687 pd=0.76 as=0.0594 ps=0.69 w=0.36 l=0.15
X3248 a_2320_16183# a_2133_15823# a_2233_15939# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.107825 ps=1.36 w=0.42 l=0.15
X3252 a_2044_15279# temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref.TE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X3255 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref.Z temp1.dac.parallel_cells\[1\].vdac_batch.einvp_batch\[0\].pupd.A a_5796_15823# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X3262 vssd1 temp1.capload\[7\].cap.TE a_6559_14735# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X3263 a_2104_26677# _114_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X3267 vssd1 del1.delay_chain\[0\].inv2.A del1.delay_chain\[1\].inv1.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X3268 a_7636_17999# a_7387_17999# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X3269 vssd1 temp1.dac.parallel_cells\[1\].vdac_batch.einvp_batch\[0\].pupd.TE a_5547_15823# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X3273 vssd1 _079_.C a_2421_13109# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X3277 a_2047_22717# _066_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1013 ps=0.99 w=0.42 l=0.15
X3283 del2.delay_chain\[0\].inv1.A a_2879_9839# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X3285 a_6735_16911# temp1.dcdc.Z temp1.capload\[8\].cap.Z vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.27 ps=2.54 w=1 l=0.15
X3288 a_4668_17143# temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[1\].pupd.TE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
R16 temp1.capload\[3\].cap_12.LO vssd1 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X3293 a_5724_17455# temp1.dac.parallel_cells\[1\].vdac_batch.einvp_batch\[1\].vref.TE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X3299 vccd1 clkbuf_1_1__f_io_in[0].A a_1674_2767# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3300 _111_.A a_4558_1653# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1625 ps=1.325 w=1 l=0.15
X3305 a_2007_11690# _063_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X3312 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[4\].pupd.A _051_.B1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3315 vccd1 del1.delay_chain\[3\].inv2.A _048_.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.25
X3317 temp1.capload\[9\].cap.Z temp1.dcdc.Z a_7636_17999# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X3333 vssd1 _053_.A1 a_1959_9615# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3334 vccd1 a_6784_17143# a_6735_16911# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1825 ps=1.365 w=1 l=0.15
X3335 a_4776_14165# _110_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.101875 ps=0.99 w=0.42 l=0.15
X3336 a_1860_14191# temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[4\].pupd.TE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X3338 a_1757_3311# a_1591_3311# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X3341 vssd1 _046_.A a_3983_18543# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X3343 vccd1 io_in[3] a_1591_7663# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X3349 a_21068_15823# a_20819_15823# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
R17 vccd1 temp1.capload\[4\].cap_13.HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X3351 vssd1 _093_.CLK a_1591_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X3352 io_out[2] a_1736_23413# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X3359 a_4157_13149# _083_.C_N vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X3369 a_1766_2223# io_in[0] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=0.15
X3373 vssd1 _111_.A a_4771_20719# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3378 del1.delay_chain\[0\].inv2.A _111_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X3379 a_4422_1501# a_3983_1135# a_4337_1135# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X3381 a_4307_12167# _051_.B1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.10025 ps=0.985 w=0.42 l=0.15
X3382 del1.delay_chain\[2\].inv1.A del1.delay_chain\[1\].inv1.Y vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X3395 vccd1 a_1674_1135# _095_.CLK vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X3396 vccd1 a_5015_1403# _110_.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3398 vssd1 a_1674_1135# _095_.CLK vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3407 vccd1 del1.delay_chain\[3\].inv2.A _048_.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.25
X3410 vssd1 temp1.dac.parallel_cells\[1\].vdac_batch.einvp_batch\[0\].pupd.TE a_5547_15279# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X3411 a_4387_1679# a_3523_1685# a_4130_1653# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X3414 del1.delay_chain\[3\].inv2.A del1.delay_chain\[2\].inv2.Y vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X3416 a_2392_16183# _085_.A1 a_2320_16183# vssd1 sky130_fd_pr__nfet_01v8 ad=0.05355 pd=0.675 as=0.0441 ps=0.63 w=0.42 l=0.15
X3417 _061_.B1_N a_1591_3855# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X3425 vssd1 temp1.capload\[4\].cap_13.LO a_7379_18543# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.235625 ps=1.375 w=0.65 l=0.15
X3432 a_2835_25236# _044_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X3434 a_7011_16617# temp1.dcdc.Z temp1.capload\[3\].cap.Z vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.27 ps=2.54 w=1 l=0.15
X3435 clkbuf_1_1__f_io_in[0].A a_1766_2223# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3437 vssd1 a_1919_22325# _067_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.169 ps=1.82 w=0.65 l=0.15
X3438 a_4516_2057# a_3523_1685# a_4387_1679# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0657 ps=0.725 w=0.36 l=0.15
X3441 a_4548_1135# a_4149_1135# a_4422_1501# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X3442 vssd1 _111_.A a_4433_21583# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3450 _115_.A a_2623_1653# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3458 vccd1 a_7980_13879# a_7931_13647# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1825 ps=1.365 w=1 l=0.15
X3460 a_4130_1653# a_3971_1679# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.1493 ps=1.22 w=0.64 l=0.15
X3474 a_4776_14165# a_4627_14191# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3475 a_4387_1679# a_3689_1685# a_4130_1653# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0657 pd=0.725 as=0.0989 ps=0.995 w=0.36 l=0.15
X3478 vssd1 _061_.B1_N a_2956_11445# vssd1 sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
X3486 a_5722_14191# _075_.A2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.095875 pd=0.945 as=0.17225 ps=1.83 w=0.65 l=0.15
X3488 _069_.A a_1715_8779# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1118 ps=1.04 w=0.65 l=0.15
X3492 a_2141_14851# _080_.A1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.074375 pd=0.815 as=0.0567 ps=0.69 w=0.42 l=0.15
X3493 vssd1 a_4590_1247# a_4548_1135# vssd1 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X3495 vccd1 a_1674_2767# _093_.CLK vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X3497 a_2406_10383# _066_.A_N a_2103_10615# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1525 pd=1.305 as=0.195 ps=1.39 w=1 l=0.15
X3499 input7.X a_1591_13647# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X3505 a_4208_19319# temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref.Z vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X3508 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref.Z temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref.Z a_5724_17455# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X3527 a_2011_10901# _111_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.2279 ps=1.74 w=0.42 l=0.15
X3532 vccd1 a_2828_20407# a_2779_20175# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1825 ps=1.365 w=1 l=0.15
X3535 a_2840_26677# _115_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X3536 vccd1 a_1828_23957# io_out[3] vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.135 ps=1.27 w=1 l=0.15
X3541 a_4418_16367# _090_.A2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.104 ps=0.97 w=0.65 l=0.15
X3549 a_3698_21583# _051_.A2 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.095875 pd=0.945 as=0.17225 ps=1.83 w=0.65 l=0.15
X3550 vccd1 a_6239_18708# temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[1\].pupd.TE vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X3551 vssd1 _066_.A_N a_2321_10703# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10075 ps=0.96 w=0.65 l=0.15
X3558 vccd1 _057_.A1 a_2222_12559# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1525 ps=1.305 w=1 l=0.15
X3562 vssd1 _095_.CLK a_3523_1685# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X3566 vccd1 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref.TE a_1683_16367# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X3574 vssd1 temp1.capload\[9\].cap.TE a_7387_17999# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
R18 temp1.capload\[0\].cap_9.HI vccd1 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X3584 a_1945_1679# _063_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X3587 _044_.A a_2327_21807# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X3588 del1.delay_chain\[1\].inv1.Y del1.delay_chain\[1\].inv1.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X3589 a_4171_18543# _111_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.2535 pd=2.08 as=0.08775 ps=0.92 w=0.65 l=0.15
X3596 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref.Z temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[4\].pupd.A a_2872_15279# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X3598 a_4413_20719# _046_.A _066_.A_N vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3612 temp1.capload\[6\].cap.Z temp1.dcdc.Z a_7012_16143# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X3613 a_4337_1135# _061_.X vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X3616 a_4215_11703# a_4487_11561# a_4445_11587# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X3629 a_4307_12167# a_4579_11995# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3634 vccd1 io_in[2] a_1591_6031# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X3640 vssd1 a_2104_25045# io_out[4] vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X3643 a_1828_23957# _112_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X3644 vccd1 temp1.capload\[6\].cap_15.LO a_6835_15823# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X3647 _112_.A _048_.B vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3651 a_1736_23413# _111_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X3658 _095_.CLK a_1674_1135# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3659 a_4619_16911# temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[1\].pupd.A temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref.Z vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.27 ps=2.54 w=1 l=0.15
X3662 vccd1 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[4\].pupd.TE a_3063_15823# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X3664 vccd1 a_3656_20407# a_3607_20175# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1825 ps=1.365 w=1 l=0.15
X3670 vccd1 a_4558_1653# _111_.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X3675 a_1674_1135# clkbuf_1_1__f_io_in[0].A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3676 vssd1 io_in[3] a_1591_7663# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X3686 vssd1 a_1766_2223# clkbuf_1_1__f_io_in[0].A vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3693 a_2593_16413# _091_.A_N vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1087 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X3696 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref.TE _109_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X3703 _093_.CLK a_1674_2767# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3706 a_7060_16519# temp1.capload\[3\].cap_12.LO vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.32075 ps=1.685 w=0.42 l=0.15
X3718 vssd1 _109_.A temp1.dac.parallel_cells\[0\].vdac_batch.einvp_batch\[0\].vref.TE vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X3719 a_4442_12265# _051_.B1 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.14825 ps=1.34 w=0.42 l=0.15
X3720 vccd1 a_1766_2223# clkbuf_1_1__f_io_in[0].A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3721 vssd1 io_in[0] a_1766_2223# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3726 vccd1 a_4031_13866# input6.X vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X3727 a_6551_15279# temp1.dcdc.Z temp1.capload\[0\].cap.Z vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.1755 ps=1.84 w=0.65 l=0.15
X3729 a_3339_13763# _110_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.14825 ps=1.34 w=0.42 l=0.15
X3730 _061_.X a_2890_11471# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X3732 vssd1 io_in[2] a_1591_6031# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X3734 a_3339_12879# _066_.A_N vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.08775 ps=0.92 w=0.65 l=0.15
X3738 vssd1 _109_.A temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref.TE vssd1 sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.091 ps=0.93 w=0.65 l=0.15
X3746 a_2828_20407# temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref.TE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X3751 vssd1 temp1.capload\[8\].cap.TE a_6735_17231# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.235625 ps=1.375 w=0.65 l=0.15
X3758 a_2835_25236# _044_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X3761 io_out[3] a_1828_23957# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X3763 a_2041_14735# _109_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1087 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X3765 vssd1 _051_.B1 temp1.dac.parallel_cells\[1\].vdac_batch.einvp_batch\[0\].pupd.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3766 a_4771_20719# _111_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3773 vccd1 _079_.B a_4579_11995# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X3776 vccd1 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref.TE a_2327_19087# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X3778 vccd1 temp1.dcdc.Z temp1.inv2.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X3781 vccd1 a_5015_1403# a_4931_1501# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X3782 a_6784_17143# temp1.capload\[8\].cap.TE vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.32075 ps=1.685 w=0.42 l=0.15
X3785 vccd1 _110_.A a_2392_13763# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X3792 a_1828_23957# _112_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
X3793 vssd1 a_1674_2767# _093_.CLK vssd1 sky130_fd_pr__nfet_01v8 ad=0.05775 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X3796 vssd1 _115_.A _066_.A_N vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3797 a_3012_17143# temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[3\].vref.TE vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.32075 ps=1.685 w=0.42 l=0.15
X3822 vccd1 _090_.A2 a_3984_16617# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3823 a_4064_1679# a_3523_1685# a_3971_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.06615 ps=0.735 w=0.42 l=0.15
X3825 _066_.A_N _046_.A a_4413_20719# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3829 _072_.C_N a_2132_9295# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.3275 ps=1.655 w=1 l=0.15
X3832 vssd1 _085_.A2 a_2392_16183# vssd1 sky130_fd_pr__nfet_01v8 ad=0.122275 pd=1.08 as=0.05355 ps=0.675 w=0.42 l=0.15
X3836 a_2818_11471# _115_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.28 ps=2.56 w=1 l=0.15
X3837 a_4771_20719# _048_.A a_4413_20719# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3838 vccd1 _090_.A2 a_3984_16617# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.145 pd=1.29 as=0.155 ps=1.31 w=1 l=0.15
X3846 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref.Z temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref.Z a_2044_18319# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X3849 a_3971_1679# a_3523_1685# a_3877_1679# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X3865 a_2872_15279# temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[4\].pupd.TE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X3866 del2.delay_chain\[0\].inv2.A del2.delay_chain\[0\].inv1.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X3870 a_1768_17231# temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref.TE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X3871 a_3984_16617# _090_.A2 vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X3884 a_2132_9295# _048_.B a_1959_9615# vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X3885 a_1959_10205# _061_.B1_N vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X3888 a_7012_16143# temp1.capload\[6\].cap_15.LO vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
R19 temp1.capload\[4\].cap_13.LO vssd1 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X3897 a_3240_16143# temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[4\].pupd.TE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X3901 vssd1 a_6239_18708# temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[1\].pupd.TE vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X3903 a_7931_13647# temp1.dac.parallel_cells\[0\].vdac_batch.einvp_batch\[0\].pupd.A temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref.Z vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.27 ps=2.54 w=1 l=0.15
X3907 vssd1 _110_.A a_2421_13109# vssd1 sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X3908 vssd1 a_3983_10927# _109_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3910 a_2095_22657# _066_.A_N vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0714 ps=0.76 w=0.42 l=0.15
X3911 _048_.A del1.delay_chain\[3\].inv2.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.25
X3915 vssd1 a_1766_2223# clkbuf_1_1__f_io_in[0].A vssd1 sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
R20 temp1.capload\[8\].cap_17.HI vccd1 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X3920 a_7980_13879# temp1.dac.parallel_cells\[0\].vdac_batch.einvp_batch\[0\].pupd.TE vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.32075 ps=1.685 w=0.42 l=0.15
X3924 vssd1 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[4\].pupd.TE a_3063_17455# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X3925 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref.TE _109_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X3941 vccd1 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[4\].pupd.TE a_3155_17999# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X3942 a_3840_17143# temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[3\].vref.TE vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.32075 ps=1.685 w=0.42 l=0.15
X3945 a_2581_2057# a_1591_1685# a_2455_1679# vssd1 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X3947 a_1920_28853# _116_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X3952 vssd1 a_2840_26677# io_out[6] vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X3969 vssd1 a_2623_3579# a_2581_3311# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X3975 a_2987_14735# _060_.B temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[4\].pupd.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3978 a_3512_12559# _066_.A_N a_3421_12559# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.1525 ps=1.305 w=1 l=0.15
X3979 vccd1 _067_.A a_1959_27247# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X3980 del2.delay_chain\[2\].inv2.Y del2.delay_chain\[2\].inv2.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X3990 _061_.B1_N a_1591_3855# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X3997 a_2116_15529# a_1867_15279# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X3999 vccd1 a_2103_11989# _060_.B vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.3275 pd=1.655 as=0.28 ps=2.56 w=1 l=0.15
X4000 _065_.X a_2971_10383# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X4010 vssd1 a_1674_1135# _095_.CLK vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4016 vssd1 _111_.A a_4771_20719# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4018 _048_.A del1.delay_chain\[3\].inv2.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.25
X4023 a_4527_18319# temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[1\].pupd.A temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref.Z vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.1755 ps=1.84 w=0.65 l=0.15
X4032 vccd1 a_1674_1135# _095_.CLK vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4033 vssd1 clkbuf_1_1__f_io_in[0].A a_1674_1135# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4039 a_4031_13866# io_in[6] vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X4040 clkbuf_1_1__f_io_in[0].A a_1766_2223# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4042 vssd1 _079_.B a_3204_13879# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X4043 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref.Z temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref.Z a_2116_15529# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X4054 vssd1 a_1674_2767# _093_.CLK vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4055 a_2011_10901# a_2187_10901# a_2139_10927# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0504 ps=0.66 w=0.42 l=0.15
X4056 a_4433_21583# _048_.A _046_.B vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4058 vccd1 _090_.A1 a_3984_16617# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4061 temp1.dac.parallel_cells\[0\].vdac_batch.einvp_batch\[0\].pupd.TE a_6559_13647# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X4067 clkbuf_1_1__f_io_in[0].A a_1766_2223# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4073 vccd1 a_7428_17607# a_7379_17705# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1825 ps=1.365 w=1 l=0.15
X4075 vssd1 _068_.B a_1801_8779# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X4087 vssd1 a_5271_14743# _051_.B1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X4088 a_4259_12879# _066_.A_N vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10725 ps=0.98 w=0.65 l=0.15
X4089 _110_.A a_5015_1403# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4093 vssd1 _109_.A temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[3\].vref.TE vssd1 sky130_fd_pr__nfet_01v8 ad=0.26 pd=2.1 as=0.08775 ps=0.92 w=0.65 l=0.15
X4094 vssd1 _079_.C a_2238_13763# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X4096 a_1768_13103# temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[4\].pupd.TE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X4098 a_7932_16367# temp1.capload\[2\].cap.TE vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.097 ps=0.975 w=0.65 l=0.15
X4103 a_3331_19087# temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[4\].pupd.A temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref.Z vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.27 ps=2.54 w=1 l=0.15
X4107 _085_.A1 a_4263_13109# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0.14825 ps=1.34 w=1 l=0.15
X4109 _048_.B a_3983_18543# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4111 vssd1 a_2103_10615# _079_.B vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X4114 vssd1 temp1.capload\[1\].cap_10.LO a_8299_18319# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.235625 ps=1.375 w=0.65 l=0.15
X4116 a_1674_1135# clkbuf_1_1__f_io_in[0].A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=0.15
X4117 _113_.A _046_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4120 a_3312_15823# a_3063_15823# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
R21 temp1.capload\[1\].cap_10.HI vccd1 sky130_fd_pr__res_generic_po w=0.48 l=0.045
X4127 vccd1 _048_.B _079_.C vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.182 pd=1.92 as=0.174 ps=1.39 w=0.7 l=0.15
X4129 vccd1 del1.delay_chain\[2\].inv2.A del1.delay_chain\[2\].inv2.Y vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X4130 vccd1 a_1674_2767# _093_.CLK vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4132 vccd1 _076_.X a_6559_13647# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X4133 a_2300_15095# _080_.A1 a_2228_15095# vssd1 sky130_fd_pr__nfet_01v8 ad=0.05355 pd=0.675 as=0.0441 ps=0.63 w=0.42 l=0.15
X4135 vssd1 a_4558_1653# _111_.A vssd1 sky130_fd_pr__nfet_01v8 ad=0.092625 pd=0.935 as=0.08775 ps=0.92 w=0.65 l=0.15
X4141 a_2421_13109# _083_.C_N vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X4142 vssd1 _065_.A a_2971_10383# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X4147 _093_.CLK a_1674_2767# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.05775 ps=0.695 w=0.42 l=0.15
X4158 vccd1 a_3380_19319# a_3331_19087# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1825 ps=1.365 w=1 l=0.15
X4160 a_2780_16373# a_2593_16413# a_2693_16631# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.107825 ps=1.36 w=0.42 l=0.15
X4161 temp1.dac.vdac_single.einvp_batch\[0\].pupd.TE _051_.B1 vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4162 vccd1 a_1766_2223# clkbuf_1_1__f_io_in[0].A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
R22 vssd1 temp1.capload\[6\].cap_15.LO sky130_fd_pr__res_generic_po w=0.48 l=0.045
X4173 vccd1 a_3983_10927# _109_.A vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4179 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref.Z temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[4\].pupd.A a_3312_15823# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X4184 a_3877_1679# _065_.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.74 as=0.1092 ps=1.36 w=0.42 l=0.15
X4185 _095_.CLK a_1674_1135# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
R23 vssd1 temp1.capload\[5\].cap.TE sky130_fd_pr__res_generic_po w=0.48 l=0.045
X4198 a_3435_13763# _079_.B a_3339_13763# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X4206 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[4\].pupd.A _060_.B a_2987_14735# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4210 a_2222_12559# _066_.A_N a_1919_12791# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1525 pd=1.305 as=0.195 ps=1.39 w=1 l=0.15
X4211 _075_.A2 a_3065_12021# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.14825 ps=1.34 w=1 l=0.15
X4215 a_4576_18231# temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[1\].pupd.TE vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.32075 ps=1.685 w=0.42 l=0.15
X4218 _061_.X a_2890_11471# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.18575 ps=1.415 w=1 l=0.15
X4219 vssd1 a_4776_14165# _090_.A1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.08775 ps=0.92 w=0.65 l=0.15
X4220 a_3689_1685# a_3523_1685# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4239 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref.Z temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref.Z a_1860_16367# vssd1 sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.235625 ps=1.375 w=0.65 l=0.15
X4240 vccd1 temp1.dac.parallel_cells\[1\].vdac_batch.einvp_batch\[0\].pupd.TE a_5547_15279# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1092 ps=1.36 w=0.42 l=0.15
X4241 a_6600_15431# temp1.capload\[0\].cap_9.LO vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X4248 _110_.A a_5015_1403# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4255 a_2007_11690# _063_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X4259 io_out[4] a_2104_25045# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.17225 ps=1.83 w=0.65 l=0.15
X4264 a_5447_18793# temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[1\].pupd.A temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref.Z vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.27 ps=2.54 w=1 l=0.15
X4266 vssd1 a_3204_13879# _080_.A2 vssd1 sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.182 ps=1.86 w=0.65 l=0.15
X4267 vssd1 a_2104_26677# io_out[5] vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.08775 ps=0.92 w=0.65 l=0.15
X4268 vssd1 a_2455_3677# a_2623_3579# vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4275 _087_.A a_2233_15939# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.122275 ps=1.08 w=0.65 l=0.15
X4280 _092_.A a_2693_16631# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142225 ps=1.335 w=1 l=0.15
X4281 vccd1 a_4387_1679# a_4558_1653# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.28 ps=2.56 w=1 l=0.15
X4282 vccd1 _090_.A1 a_3984_16617# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4283 a_2030_1679# a_1757_1685# a_1945_1679# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X4286 vccd1 a_4208_19319# a_4159_19087# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.32075 pd=1.685 as=0.1825 ps=1.365 w=1 l=0.15
X4288 a_5796_16617# a_5547_16367# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1825 pd=1.365 as=0.32075 ps=1.685 w=1 l=0.15
X4289 a_4341_12559# input7.X vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X4293 _093_.CLK a_1674_2767# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4299 io_out[7] a_1920_28853# vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X4300 temp1.dac.vdac_single.einvp_batch\[0\].pupd.TE _071_.C vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4301 vccd1 _093_.CLK a_1591_1685# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X4307 a_7379_18543# temp1.dcdc.Z temp1.capload\[4\].cap.Z vssd1 sky130_fd_pr__nfet_01v8 ad=0.235625 pd=1.375 as=0.1755 ps=1.84 w=0.65 l=0.15
X4308 vssd1 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref.TE a_1867_17999# vssd1 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X4325 _051_.B1 a_5271_14743# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X4327 temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[3\].vref.TE _109_.A vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10725 ps=0.98 w=0.65 l=0.15
X4331 vssd1 _067_.A a_1959_27247# vssd1 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X4332 a_2852_16373# _090_.A1 a_2780_16373# vssd1 sky130_fd_pr__nfet_01v8 ad=0.05355 pd=0.675 as=0.0441 ps=0.63 w=0.42 l=0.15
X4338 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref.Z temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref.Z a_5796_16617# vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.1825 ps=1.365 w=1 l=0.15
X4344 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[4\].pupd.TE a_5323_17973# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X4347 _095_.CLK a_1674_1135# vssd1 vssd1 sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4349 a_2932_21237# _109_.A vccd1 vccd1 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.149 ps=1.325 w=0.64 l=0.15
C0 a_4337_1135# vssd1 0.23fF $ **FLOATING
C1 a_4847_1501# vssd1 0.61fF $ **FLOATING
C2 a_5015_1403# vssd1 0.97fF $ **FLOATING
C3 a_4422_1501# vssd1 0.63fF $ **FLOATING
C4 a_4590_1247# vssd1 0.58fF $ **FLOATING
C5 a_4149_1135# vssd1 1.43fF $ **FLOATING
C6 a_3983_1135# vssd1 1.81fF $ **FLOATING
C7 a_1674_1135# vssd1 4.03fF $ **FLOATING
C8 a_3877_1679# vssd1 0.22fF $ **FLOATING
C9 a_1945_1679# vssd1 0.23fF $ **FLOATING
C10 a_4387_1679# vssd1 0.60fF $ **FLOATING
C11 a_4558_1653# vssd1 1.41fF $ **FLOATING
C12 a_3971_1679# vssd1 0.63fF $ **FLOATING
C13 a_4130_1653# vssd1 0.59fF $ **FLOATING
C14 a_3689_1685# vssd1 1.39fF $ **FLOATING
C15 a_3523_1685# vssd1 1.77fF $ **FLOATING
C16 _095_.CLK vssd1 3.46fF $ **FLOATING
C17 a_2455_1679# vssd1 0.61fF $ **FLOATING
C18 a_2623_1653# vssd1 0.97fF $ **FLOATING
C19 a_2030_1679# vssd1 0.63fF $ **FLOATING
C20 a_2198_1653# vssd1 0.58fF $ **FLOATING
C21 a_1757_1685# vssd1 1.43fF $ **FLOATING
C22 a_1591_1685# vssd1 1.81fF $ **FLOATING
C23 a_1766_2223# vssd1 4.03fF $ **FLOATING
C24 io_in[0] vssd1 2.01fF
C25 a_1674_2767# vssd1 4.03fF $ **FLOATING
C26 clkbuf_1_1__f_io_in[0].A vssd1 5.28fF $ **FLOATING
C27 a_1945_3311# vssd1 0.23fF $ **FLOATING
C28 a_2455_3677# vssd1 0.61fF $ **FLOATING
C29 a_2623_3579# vssd1 0.82fF $ **FLOATING
C30 a_2030_3677# vssd1 0.63fF $ **FLOATING
C31 a_2198_3423# vssd1 0.58fF $ **FLOATING
C32 a_1757_3311# vssd1 1.43fF $ **FLOATING
C33 a_1591_3311# vssd1 1.81fF $ **FLOATING
C34 _093_.CLK vssd1 4.20fF $ **FLOATING
C35 a_1591_3855# vssd1 0.52fF $ **FLOATING
C36 io_in[1] vssd1 1.32fF
C37 a_1591_6031# vssd1 0.52fF $ **FLOATING
C38 io_in[2] vssd1 1.38fF
C39 a_1591_7663# vssd1 0.52fF $ **FLOATING
C40 io_in[3] vssd1 1.18fF
C41 _068_.B vssd1 1.70fF $ **FLOATING
C42 a_1715_8779# vssd1 0.56fF $ **FLOATING
C43 a_1959_9615# vssd1 0.17fF $ **FLOATING
C44 io_in[4] vssd1 1.92fF
C45 a_2927_9514# vssd1 0.52fF $ **FLOATING
C46 a_2132_9295# vssd1 0.55fF $ **FLOATING
C47 _053_.A1 vssd1 1.30fF $ **FLOATING
C48 a_2879_9839# vssd1 0.52fF $ **FLOATING
C49 _069_.A vssd1 1.44fF $ **FLOATING
C50 a_2139_10205# vssd1 0.51fF $ **FLOATING
C51 a_1959_10205# vssd1 0.60fF $ **FLOATING
C52 _065_.X vssd1 4.35fF $ **FLOATING
C53 a_2321_10703# vssd1 0.17fF $ **FLOATING
C54 del2.delay_chain\[0\].inv1.A vssd1 1.28fF $ **FLOATING
C55 a_2971_10383# vssd1 0.52fF $ **FLOATING
C56 _065_.A vssd1 1.08fF $ **FLOATING
C57 _055_.A1 vssd1 1.16fF $ **FLOATING
C58 a_2103_10615# vssd1 0.55fF $ **FLOATING
C59 a_3983_10927# vssd1 1.20fF $ **FLOATING
C60 io_in[5] vssd1 2.11fF
C61 a_2927_11092# vssd1 0.52fF $ **FLOATING
C62 a_2187_10901# vssd1 0.60fF $ **FLOATING
C63 a_2011_10901# vssd1 0.51fF $ **FLOATING
C64 del2.delay_chain\[0\].inv2.A vssd1 1.45fF $ **FLOATING
C65 a_4487_11561# vssd1 0.43fF $ **FLOATING
C66 _061_.X vssd1 5.20fF $ **FLOATING
C67 _061_.B1_N vssd1 6.14fF $ **FLOATING
C68 a_2723_11791# vssd1 0.20fF $ **FLOATING
C69 _063_.X vssd1 4.65fF $ **FLOATING
C70 a_4215_11703# vssd1 0.67fF $ **FLOATING
C71 a_2890_11471# vssd1 0.65fF $ **FLOATING
C72 a_2956_11445# vssd1 0.44fF $ **FLOATING
C73 _063_.A vssd1 0.92fF $ **FLOATING
C74 a_2007_11690# vssd1 0.52fF $ **FLOATING
C75 a_2321_12015# vssd1 0.17fF $ **FLOATING
C76 a_4579_11995# vssd1 0.43fF $ **FLOATING
C77 _072_.C_N vssd1 4.27fF $ **FLOATING
C78 a_4307_12167# vssd1 0.67fF $ **FLOATING
C79 a_3065_12021# vssd1 0.66fF $ **FLOATING
C80 a_2103_11989# vssd1 0.55fF $ **FLOATING
C81 a_4259_12879# vssd1 0.18fF $ **FLOATING
C82 a_3339_12879# vssd1 0.17fF $ **FLOATING
C83 a_2137_12879# vssd1 0.17fF $ **FLOATING
C84 a_3512_12559# vssd1 0.55fF $ **FLOATING
C85 _057_.A1 vssd1 1.45fF $ **FLOATING
C86 a_1919_12791# vssd1 0.55fF $ **FLOATING
C87 a_4157_13149# vssd1 0.43fF $ **FLOATING
C88 a_4263_13109# vssd1 0.67fF $ **FLOATING
C89 _083_.C_N vssd1 2.55fF $ **FLOATING
C90 a_2421_13109# vssd1 0.66fF $ **FLOATING
C91 a_1591_13103# vssd1 0.53fF $ **FLOATING
C92 a_7980_13879# vssd1 0.53fF $ **FLOATING
C93 input6.X vssd1 1.84fF $ **FLOATING
C94 temp1.dac.parallel_cells\[0\].vdac_batch.einvp_batch\[0\].pupd.TE vssd1 1.48fF $ **FLOATING
C95 temp1.dac.parallel_cells\[0\].vdac_batch.einvp_batch\[0\].pupd.A vssd1 2.97fF $ **FLOATING
C96 a_6559_13647# vssd1 0.52fF $ **FLOATING
C97 a_5271_13647# vssd1 0.52fF $ **FLOATING
C98 io_in[6] vssd1 2.29fF
C99 a_4031_13866# vssd1 0.52fF $ **FLOATING
C100 _079_.B vssd1 4.20fF $ **FLOATING
C101 a_3204_13879# vssd1 0.66fF $ **FLOATING
C102 a_2238_13763# vssd1 0.82fF $ **FLOATING
C103 _079_.C vssd1 4.04fF $ **FLOATING
C104 input7.X vssd1 2.37fF $ **FLOATING
C105 a_1591_13647# vssd1 0.52fF $ **FLOATING
C106 io_in[7] vssd1 1.98fF
C107 a_7479_14191# vssd1 0.53fF $ **FLOATING
C108 temp1.capload\[7\].cap_16.HI vssd1 0.42fF $ **FLOATING
C109 temp1.dac.parallel_cells\[0\].vdac_batch.einvp_batch\[0\].vref.TE vssd1 1.52fF $ **FLOATING
C110 a_5639_14441# vssd1 0.24fF $ **FLOATING
C111 a_4627_14191# vssd1 0.73fF $ **FLOATING
C112 _076_.X vssd1 2.23fF $ **FLOATING
C113 _075_.A2 vssd1 2.82fF $ **FLOATING
C114 a_4776_14165# vssd1 0.72fF $ **FLOATING
C115 a_2877_14455# vssd1 0.60fF $ **FLOATING
C116 _075_.A1 vssd1 3.60fF $ **FLOATING
C117 a_2777_14237# vssd1 0.49fF $ **FLOATING
C118 a_1683_14191# vssd1 0.53fF $ **FLOATING
C119 a_4535_14735# vssd1 0.24fF $ **FLOATING
C120 a_2987_14735# vssd1 0.39fF $ **FLOATING
C121 temp1.capload\[7\].cap.Z vssd1 0.29fF $ **FLOATING
C122 a_6559_14735# vssd1 0.53fF $ **FLOATING
C123 _081_.X vssd1 2.21fF $ **FLOATING
C124 temp1.capload\[7\].cap.TE vssd1 1.28fF $ **FLOATING
C125 a_5271_14743# vssd1 0.65fF $ **FLOATING
C126 _071_.C vssd1 4.91fF $ **FLOATING
C127 _060_.B vssd1 3.94fF $ **FLOATING
C128 a_2141_14851# vssd1 0.60fF $ **FLOATING
C129 _080_.A2 vssd1 2.68fF $ **FLOATING
C130 _080_.A1 vssd1 3.69fF $ **FLOATING
C131 a_2041_14735# vssd1 0.49fF $ **FLOATING
C132 temp1.capload\[0\].cap_9.HI vssd1 0.42fF $ **FLOATING
C133 temp1.capload\[8\].cap_17.HI vssd1 0.42fF $ **FLOATING
C134 temp1.capload\[0\].cap.Z vssd1 0.29fF $ **FLOATING
C135 a_4443_15529# vssd1 0.44fF $ **FLOATING
C136 temp1.capload\[0\].cap_9.LO vssd1 1.51fF $ **FLOATING
C137 a_6600_15431# vssd1 0.53fF $ **FLOATING
C138 a_5547_15279# vssd1 0.53fF $ **FLOATING
C139 a_2695_15279# vssd1 0.53fF $ **FLOATING
C140 a_1867_15279# vssd1 0.53fF $ **FLOATING
C141 a_20819_15823# vssd1 0.53fF $ **FLOATING
C142 temp1.dac.vdac_single.einvp_batch\[0\].pupd.TE vssd1 9.00fF $ **FLOATING
C143 temp1.capload\[2\].cap_11.HI vssd1 0.42fF $ **FLOATING
C144 temp1.capload\[6\].cap.Z vssd1 0.29fF $ **FLOATING
C145 a_6835_15823# vssd1 0.53fF $ **FLOATING
C146 a_5547_15823# vssd1 0.53fF $ **FLOATING
C147 a_4535_15823# vssd1 0.53fF $ **FLOATING
C148 a_3063_15823# vssd1 0.53fF $ **FLOATING
C149 temp1.dac.parallel_cells\[1\].vdac_batch.einvp_batch\[0\].pupd.A vssd1 2.76fF $ **FLOATING
C150 temp1.dac.parallel_cells\[1\].vdac_batch.einvp_batch\[0\].pupd.TE vssd1 2.33fF $ **FLOATING
C151 del2.delay_chain\[1\].inv1.A vssd1 2.80fF $ **FLOATING
C152 a_2233_15939# vssd1 0.60fF $ **FLOATING
C153 _085_.A2 vssd1 3.28fF $ **FLOATING
C154 _085_.A1 vssd1 3.21fF $ **FLOATING
C155 a_2133_15823# vssd1 0.49fF $ **FLOATING
C156 temp1.dac.vdac_single.einvp_batch\[0\].pupd_20.LO vssd1 0.48fF $ **FLOATING
C157 temp1.dac.vdac_single.einvp_batch\[0\].pupd_20.HI vssd1 1.06fF $ **FLOATING
C158 temp1.capload\[2\].cap.Z vssd1 0.29fF $ **FLOATING
C159 a_4418_16367# vssd1 0.36fF $ **FLOATING
C160 temp1.capload\[3\].cap.Z vssd1 0.29fF $ **FLOATING
C161 a_3984_16617# vssd1 0.71fF $ **FLOATING
C162 a_9135_16367# vssd1 0.53fF $ **FLOATING
C163 a_7755_16367# vssd1 0.53fF $ **FLOATING
C164 temp1.capload\[2\].cap.TE vssd1 1.38fF $ **FLOATING
C165 a_7060_16519# vssd1 0.53fF $ **FLOATING
C166 a_5547_16367# vssd1 0.53fF $ **FLOATING
C167 _090_.A2 vssd1 4.53fF $ **FLOATING
C168 a_2693_16631# vssd1 0.60fF $ **FLOATING
C169 _090_.A1 vssd1 3.39fF $ **FLOATING
C170 a_2593_16413# vssd1 0.49fF $ **FLOATING
C171 _091_.A_N vssd1 7.28fF $ **FLOATING
C172 a_1683_16367# vssd1 0.53fF $ **FLOATING
C173 temp1.dac.vdac_single.einvp_batch\[0\].vref_19.LO vssd1 1.52fF $ **FLOATING
C174 temp1.dac.vdac_single.einvp_batch\[0\].vref_19.HI vssd1 0.42fF $ **FLOATING
C175 temp1.capload\[3\].cap_12.HI vssd1 0.42fF $ **FLOATING
C176 temp1.capload\[3\].cap_12.LO vssd1 1.36fF $ **FLOATING
C177 a_6784_17143# vssd1 0.53fF $ **FLOATING
C178 temp1.capload\[8\].cap.Z vssd1 0.29fF $ **FLOATING
C179 a_5547_16911# vssd1 0.53fF $ **FLOATING
C180 a_4668_17143# vssd1 0.53fF $ **FLOATING
C181 a_3840_17143# vssd1 0.53fF $ **FLOATING
C182 a_3012_17143# vssd1 0.53fF $ **FLOATING
C183 a_1591_16911# vssd1 0.53fF $ **FLOATING
C184 temp1.capload\[8\].cap.TE vssd1 1.83fF $ **FLOATING
C185 temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[3\].vref.TE vssd1 4.60fF $ **FLOATING
C186 temp1.capload\[5\].cap_14.HI vssd1 0.42fF $ **FLOATING
C187 temp1.capload\[5\].cap.Z vssd1 0.29fF $ **FLOATING
C188 temp1.capload\[5\].cap.TE vssd1 1.24fF $ **FLOATING
C189 a_7428_17607# vssd1 0.53fF $ **FLOATING
C190 temp1.capload\[6\].cap_15.LO vssd1 1.76fF $ **FLOATING
C191 temp1.capload\[6\].cap_15.HI vssd1 0.42fF $ **FLOATING
C192 a_5547_17455# vssd1 0.53fF $ **FLOATING
C193 temp1.dac.parallel_cells\[1\].vdac_batch.einvp_batch\[1\].vref.TE vssd1 2.90fF $ **FLOATING
C194 a_4535_17455# vssd1 0.53fF $ **FLOATING
C195 a_3063_17455# vssd1 0.53fF $ **FLOATING
C196 a_1867_17455# vssd1 0.53fF $ **FLOATING
C197 a_8348_18231# vssd1 0.53fF $ **FLOATING
C198 temp1.capload\[1\].cap.Z vssd1 0.29fF $ **FLOATING
C199 temp1.capload\[9\].cap.Z vssd1 0.29fF $ **FLOATING
C200 a_7387_17999# vssd1 0.53fF $ **FLOATING
C201 temp1.capload\[9\].cap.TE vssd1 1.24fF $ **FLOATING
C202 temp1.capload\[9\].cap_18.HI vssd1 0.42fF $ **FLOATING
C203 a_4576_18231# vssd1 0.53fF $ **FLOATING
C204 a_3155_17999# vssd1 0.53fF $ **FLOATING
C205 a_1867_17999# vssd1 0.53fF $ **FLOATING
C206 _092_.A vssd1 2.28fF $ **FLOATING
C207 a_5323_17973# vssd1 0.70fF $ **FLOATING
C208 temp1.capload\[1\].cap_10.LO vssd1 1.45fF $ **FLOATING
C209 temp1.capload\[1\].cap_10.HI vssd1 0.42fF $ **FLOATING
C210 a_4171_18543# vssd1 0.52fF $ **FLOATING
C211 temp1.capload\[4\].cap.Z vssd1 0.29fF $ **FLOATING
C212 a_7428_18695# vssd1 0.53fF $ **FLOATING
C213 _087_.A vssd1 3.50fF $ **FLOATING
C214 a_6239_18708# vssd1 0.52fF $ **FLOATING
C215 temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[1\].pupd.TE vssd1 3.99fF $ **FLOATING
C216 a_5496_18695# vssd1 0.53fF $ **FLOATING
C217 temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[1\].pupd.A vssd1 5.34fF $ **FLOATING
C218 a_3983_18543# vssd1 1.14fF $ **FLOATING
C219 a_3063_18543# vssd1 0.53fF $ **FLOATING
C220 temp1.capload\[4\].cap_13.LO vssd1 1.32fF $ **FLOATING
C221 temp1.capload\[4\].cap_13.HI vssd1 0.42fF $ **FLOATING
C222 a_4208_19319# vssd1 0.53fF $ **FLOATING
C223 a_3380_19319# vssd1 0.53fF $ **FLOATING
C224 a_2327_19087# vssd1 0.53fF $ **FLOATING
C225 temp1.dcdc.Z vssd1 8.91fF $ **FLOATING
C226 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[4\].pupd.TE vssd1 9.18fF $ **FLOATING
C227 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[4\].pupd.A vssd1 6.65fF $ **FLOATING
C228 del1.delay_chain\[3\].inv2.A vssd1 1.73fF $ **FLOATING
C229 a_3656_20407# vssd1 0.53fF $ **FLOATING
C230 a_2828_20407# vssd1 0.53fF $ **FLOATING
C231 del1.delay_chain\[2\].inv1.A vssd1 2.21fF $ **FLOATING
C232 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref.TE vssd1 9.21fF $ **FLOATING
C233 temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref.Z vssd1 35.66fF $ **FLOATING
C234 a_4771_20719# vssd1 0.43fF $ **FLOATING
C235 a_4413_20719# vssd1 0.31fF $ **FLOATING
C236 a_3983_20969# vssd1 1.23fF $ **FLOATING
C237 del1.delay_chain\[2\].inv2.Y vssd1 1.23fF $ **FLOATING
C238 del1.delay_chain\[0\].inv2.A vssd1 1.22fF $ **FLOATING
C239 del1.delay_chain\[2\].inv2.A vssd1 1.89fF $ **FLOATING
C240 a_3615_21263# vssd1 0.24fF $ **FLOATING
C241 _051_.Y vssd1 1.60fF $ **FLOATING
C242 io_out[0] vssd1 2.97fF
C243 del1.delay_chain\[1\].inv1.Y vssd1 1.68fF $ **FLOATING
C244 _051_.B1 vssd1 12.54fF $ **FLOATING
C245 _051_.A2 vssd1 0.97fF $ **FLOATING
C246 _109_.A vssd1 13.65fF $ **FLOATING
C247 a_2932_21237# vssd1 0.65fF $ **FLOATING
C248 del1.delay_chain\[1\].inv1.A vssd1 0.99fF $ **FLOATING
C249 del2.delay_chain\[1\].inv2.Y vssd1 3.92fF $ **FLOATING
C250 temp1.inv2.A vssd1 1.97fF $ **FLOATING
C251 del2.delay_chain\[1\].inv2.A vssd1 3.20fF $ **FLOATING
C252 a_2327_21807# vssd1 0.62fF $ **FLOATING
C253 _110_.A vssd1 14.85fF $ **FLOATING
C254 io_out[1] vssd1 1.84fF
C255 a_1644_21781# vssd1 0.65fF $ **FLOATING
C256 del2.delay_chain\[3\].inv2.A vssd1 2.47fF $ **FLOATING
C257 _066_.A_N vssd1 11.51fF $ **FLOATING
C258 a_2095_22657# vssd1 0.60fF $ **FLOATING
C259 _066_.B vssd1 1.77fF $ **FLOATING
C260 a_1919_22325# vssd1 0.51fF $ **FLOATING
C261 del2.delay_chain\[2\].inv2.Y vssd1 1.66fF $ **FLOATING
C262 _048_.A vssd1 10.37fF $ **FLOATING
C263 _048_.B vssd1 11.32fF $ **FLOATING
C264 del2.delay_chain\[2\].inv2.A vssd1 4.90fF $ **FLOATING
C265 io_out[2] vssd1 1.72fF
C266 _046_.B vssd1 2.53fF $ **FLOATING
C267 _046_.A vssd1 6.24fF $ **FLOATING
C268 _111_.A vssd1 17.11fF $ **FLOATING
C269 a_1736_23413# vssd1 0.65fF $ **FLOATING
C270 _112_.A vssd1 1.30fF $ **FLOATING
C271 io_out[3] vssd1 1.26fF
C272 a_1828_23957# vssd1 0.65fF $ **FLOATING
C273 _044_.A vssd1 2.13fF $ **FLOATING
C274 a_2835_25236# vssd1 0.52fF $ **FLOATING
C275 _113_.A vssd1 1.40fF $ **FLOATING
C276 io_out[4] vssd1 1.61fF
C277 a_2104_25045# vssd1 0.65fF $ **FLOATING
C278 io_out[6] vssd1 2.88fF
C279 io_out[5] vssd1 2.33fF
C280 _115_.A vssd1 13.38fF $ **FLOATING
C281 a_2840_26677# vssd1 0.65fF $ **FLOATING
C282 _114_.A vssd1 1.50fF $ **FLOATING
C283 a_2104_26677# vssd1 0.65fF $ **FLOATING
C284 a_1959_27247# vssd1 0.52fF $ **FLOATING
C285 _067_.A vssd1 2.55fF $ **FLOATING
C286 io_out[7] vssd1 3.15fF
C287 _116_.A vssd1 1.32fF $ **FLOATING
C288 a_1920_28853# vssd1 0.65fF $ **FLOATING
C289 vccd1 vssd1 4386.08fF
.ends
